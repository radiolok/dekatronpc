module DekatronPulseAllow(
    input wire CarryLow,
    input wire CarryHigh,
    input wire Dec,//High if Dec
    //Input pulses:
    input wire [1:0] PulsesIn,
    //Output pulses:
    output wire [1:0] PulsesOut
);
endmodule
