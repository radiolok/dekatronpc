module pi(Address, Data);

parameter portSize = 12;
parameter dataSize = 4;

/* verilator lint_off UNUSEDSIGNAL */
input logic [portSize-1:0] Address;
/* verilator lint_on UNUSEDSIGNAL */
output logic [dataSize-1:0] Data;

always_comb
/* verilator lint_off WIDTHEXPAND */
  case(Address)
    12'b0000: Data = {4'b0010}; //+
    12'b0001: Data = {4'b0010}; //+
    12'b0010: Data = {4'b0010}; //+
    12'b0011: Data = {4'b0010}; //+
    12'b0100: Data = {4'b0110}; //[
    12'b0101: Data = {4'b0101}; //<
    12'b0110: Data = {4'b0010}; //+
    12'b0111: Data = {4'b0100}; //>
    12'b1000: Data = {4'b0100}; //>
    12'b1001: Data = {4'b0100}; //>
    12'b00010000: Data = {4'b0100}; //>
    12'b00010001: Data = {4'b0100}; //>
    12'b00010010: Data = {4'b0100}; //>
    12'b00010011: Data = {4'b0100}; //>
    12'b00010100: Data = {4'b0100}; //>
    12'b00010101: Data = {4'b0010}; //+
    12'b00010110: Data = {4'b0010}; //+
    12'b00010111: Data = {4'b0010}; //+
    12'b00011000: Data = {4'b0010}; //+
    12'b00011001: Data = {4'b0010}; //+
    12'b00100000: Data = {4'b0010}; //+
    12'b00100001: Data = {4'b0010}; //+
    12'b00100010: Data = {4'b0010}; //+
    12'b00100011: Data = {4'b0010}; //+
    12'b00100100: Data = {4'b0010}; //+
    12'b00100101: Data = {4'b0101}; //<
    12'b00100110: Data = {4'b0101}; //<
    12'b00100111: Data = {4'b0101}; //<
    12'b00101000: Data = {4'b0101}; //<
    12'b00101001: Data = {4'b0101}; //<
    12'b00110000: Data = {4'b0101}; //<
    12'b00110001: Data = {4'b0101}; //<
    12'b00110010: Data = {4'b0011}; //-
    12'b00110011: Data = {4'b0111}; //]
    12'b00110100: Data = {4'b0100}; //>
    12'b00110101: Data = {4'b0010}; //+
    12'b00110110: Data = {4'b0010}; //+
    12'b00110111: Data = {4'b0010}; //+
    12'b00111000: Data = {4'b0010}; //+
    12'b00111001: Data = {4'b0010}; //+
    12'b01000000: Data = {4'b0110}; //[
    12'b01000001: Data = {4'b0101}; //<
    12'b01000010: Data = {4'b0010}; //+
    12'b01000011: Data = {4'b0010}; //+
    12'b01000100: Data = {4'b0010}; //+
    12'b01000101: Data = {4'b0010}; //+
    12'b01000110: Data = {4'b0010}; //+
    12'b01000111: Data = {4'b0010}; //+
    12'b01001000: Data = {4'b0010}; //+
    12'b01001001: Data = {4'b0010}; //+
    12'b01010000: Data = {4'b0010}; //+
    12'b01010001: Data = {4'b0100}; //>
    12'b01010010: Data = {4'b0011}; //-
    12'b01010011: Data = {4'b0111}; //]
    12'b01010100: Data = {4'b0010}; //+
    12'b01010101: Data = {4'b0100}; //>
    12'b01010110: Data = {4'b0100}; //>
    12'b01010111: Data = {4'b0100}; //>
    12'b01011000: Data = {4'b0100}; //>
    12'b01011001: Data = {4'b0100}; //>
    12'b01100000: Data = {4'b0100}; //>
    12'b01100001: Data = {4'b0010}; //+
    12'b01100010: Data = {4'b0110}; //[
    12'b01100011: Data = {4'b0101}; //<
    12'b01100100: Data = {4'b0101}; //<
    12'b01100101: Data = {4'b0010}; //+
    12'b01100110: Data = {4'b0010}; //+
    12'b01100111: Data = {4'b0010}; //+
    12'b01101000: Data = {4'b0110}; //[
    12'b01101001: Data = {4'b0100}; //>
    12'b01110000: Data = {4'b0100}; //>
    12'b01110001: Data = {4'b0110}; //[
    12'b01110010: Data = {4'b0011}; //-
    12'b01110011: Data = {4'b0101}; //<
    12'b01110100: Data = {4'b0111}; //]
    12'b01110101: Data = {4'b0101}; //<
    12'b01110110: Data = {4'b0110}; //[
    12'b01110111: Data = {4'b0100}; //>
    12'b01111000: Data = {4'b0111}; //]
    12'b01111001: Data = {4'b0101}; //<
    12'b10000000: Data = {4'b0011}; //-
    12'b10000001: Data = {4'b0111}; //]
    12'b10000010: Data = {4'b0100}; //>
    12'b10000011: Data = {4'b0100}; //>
    12'b10000100: Data = {4'b0110}; //[
    12'b10000101: Data = {4'b0100}; //>
    12'b10000110: Data = {4'b0010}; //+
    12'b10000111: Data = {4'b0100}; //>
    12'b10001000: Data = {4'b0111}; //]
    12'b10001001: Data = {4'b0101}; //<
    12'b10010000: Data = {4'b0110}; //[
    12'b10010001: Data = {4'b0101}; //<
    12'b10010010: Data = {4'b0111}; //]
    12'b10010011: Data = {4'b0100}; //>
    12'b10010100: Data = {4'b0111}; //]
    12'b10010101: Data = {4'b0100}; //>
    12'b10010110: Data = {4'b0110}; //[
    12'b10010111: Data = {4'b0110}; //[
    12'b10011000: Data = {4'b0011}; //-
    12'b10011001: Data = {4'b0100}; //>
    12'b000100000000: Data = {4'b0100}; //>
    12'b000100000001: Data = {4'b0100}; //>
    12'b000100000010: Data = {4'b0100}; //>
    12'b000100000011: Data = {4'b0010}; //+
    12'b000100000100: Data = {4'b0101}; //<
    12'b000100000101: Data = {4'b0101}; //<
    12'b000100000110: Data = {4'b0101}; //<
    12'b000100000111: Data = {4'b0101}; //<
    12'b000100001000: Data = {4'b0111}; //]
    12'b000100001001: Data = {4'b0100}; //>
    12'b000100010000: Data = {4'b0100}; //>
    12'b000100010001: Data = {4'b0100}; //>
    12'b000100010010: Data = {4'b0010}; //+
    12'b000100010011: Data = {4'b0010}; //+
    12'b000100010100: Data = {4'b0010}; //+
    12'b000100010101: Data = {4'b0100}; //>
    12'b000100010110: Data = {4'b0011}; //-
    12'b000100010111: Data = {4'b0111}; //]
    12'b000100011000: Data = {4'b0101}; //<
    12'b000100011001: Data = {4'b0110}; //[
    12'b000100100000: Data = {4'b0101}; //<
    12'b000100100001: Data = {4'b0101}; //<
    12'b000100100010: Data = {4'b0101}; //<
    12'b000100100011: Data = {4'b0101}; //<
    12'b000100100100: Data = {4'b0111}; //]
    12'b000100100101: Data = {4'b0101}; //<
    12'b000100100110: Data = {4'b0101}; //<
    12'b000100100111: Data = {4'b0101}; //<
    12'b000100101000: Data = {4'b0101}; //<
    12'b000100101001: Data = {4'b0101}; //<
    12'b000100110000: Data = {4'b0101}; //<
    12'b000100110001: Data = {4'b0101}; //<
    12'b000100110010: Data = {4'b0101}; //<
    12'b000100110011: Data = {4'b0010}; //+
    12'b000100110100: Data = {4'b0110}; //[
    12'b000100110101: Data = {4'b0011}; //-
    12'b000100110110: Data = {4'b0100}; //>
    12'b000100110111: Data = {4'b0100}; //>
    12'b000100111000: Data = {4'b0100}; //>
    12'b000100111001: Data = {4'b0100}; //>
    12'b000101000000: Data = {4'b0100}; //>
    12'b000101000001: Data = {4'b0100}; //>
    12'b000101000010: Data = {4'b0100}; //>
    12'b000101000011: Data = {4'b0100}; //>
    12'b000101000100: Data = {4'b0100}; //>
    12'b000101000101: Data = {4'b0100}; //>
    12'b000101000110: Data = {4'b0100}; //>
    12'b000101000111: Data = {4'b0100}; //>
    12'b000101001000: Data = {4'b0110}; //[
    12'b000101001001: Data = {4'b0101}; //<
    12'b000101010000: Data = {4'b0010}; //+
    12'b000101010001: Data = {4'b0110}; //[
    12'b000101010010: Data = {4'b0011}; //-
    12'b000101010011: Data = {4'b0100}; //>
    12'b000101010100: Data = {4'b0100}; //>
    12'b000101010101: Data = {4'b0100}; //>
    12'b000101010110: Data = {4'b0100}; //>
    12'b000101010111: Data = {4'b0010}; //+
    12'b000101011000: Data = {4'b0101}; //<
    12'b000101011001: Data = {4'b0101}; //<
    12'b000101100000: Data = {4'b0101}; //<
    12'b000101100001: Data = {4'b0101}; //<
    12'b000101100010: Data = {4'b0111}; //]
    12'b000101100011: Data = {4'b0100}; //>
    12'b000101100100: Data = {4'b0100}; //>
    12'b000101100101: Data = {4'b0100}; //>
    12'b000101100110: Data = {4'b0100}; //>
    12'b000101100111: Data = {4'b0100}; //>
    12'b000101101000: Data = {4'b0111}; //]
    12'b000101101001: Data = {4'b0101}; //<
    12'b000101110000: Data = {4'b0101}; //<
    12'b000101110001: Data = {4'b0101}; //<
    12'b000101110010: Data = {4'b0101}; //<
    12'b000101110011: Data = {4'b0110}; //[
    12'b000101110100: Data = {4'b0100}; //>
    12'b000101110101: Data = {4'b0100}; //>
    12'b000101110110: Data = {4'b0100}; //>
    12'b000101110111: Data = {4'b0100}; //>
    12'b000101111000: Data = {4'b0100}; //>
    12'b000101111001: Data = {4'b0110}; //[
    12'b000110000000: Data = {4'b0101}; //<
    12'b000110000001: Data = {4'b0101}; //<
    12'b000110000010: Data = {4'b0101}; //<
    12'b000110000011: Data = {4'b0101}; //<
    12'b000110000100: Data = {4'b0010}; //+
    12'b000110000101: Data = {4'b0100}; //>
    12'b000110000110: Data = {4'b0100}; //>
    12'b000110000111: Data = {4'b0100}; //>
    12'b000110001000: Data = {4'b0100}; //>
    12'b000110001001: Data = {4'b0011}; //-
    12'b000110010000: Data = {4'b0111}; //]
    12'b000110010001: Data = {4'b0101}; //<
    12'b000110010010: Data = {4'b0101}; //<
    12'b000110010011: Data = {4'b0101}; //<
    12'b000110010100: Data = {4'b0101}; //<
    12'b000110010101: Data = {4'b0101}; //<
    12'b000110010110: Data = {4'b0011}; //-
    12'b000110010111: Data = {4'b0110}; //[
    12'b000110011000: Data = {4'b0101}; //<
    12'b000110011001: Data = {4'b0101}; //<
    12'b001000000000: Data = {4'b0010}; //+
    12'b001000000001: Data = {4'b0010}; //+
    12'b001000000010: Data = {4'b0010}; //+
    12'b001000000011: Data = {4'b0010}; //+
    12'b001000000100: Data = {4'b0010}; //+
    12'b001000000101: Data = {4'b0010}; //+
    12'b001000000110: Data = {4'b0010}; //+
    12'b001000000111: Data = {4'b0010}; //+
    12'b001000001000: Data = {4'b0010}; //+
    12'b001000001001: Data = {4'b0010}; //+
    12'b001000010000: Data = {4'b0100}; //>
    12'b001000010001: Data = {4'b0100}; //>
    12'b001000010010: Data = {4'b0011}; //-
    12'b001000010011: Data = {4'b0111}; //]
    12'b001000010100: Data = {4'b0100}; //>
    12'b001000010101: Data = {4'b0100}; //>
    12'b001000010110: Data = {4'b0100}; //>
    12'b001000010111: Data = {4'b0110}; //[
    12'b001000011000: Data = {4'b0101}; //<
    12'b001000011001: Data = {4'b0101}; //<
    12'b001000100000: Data = {4'b0110}; //[
    12'b001000100001: Data = {4'b0101}; //<
    12'b001000100010: Data = {4'b0010}; //+
    12'b001000100011: Data = {4'b0101}; //<
    12'b001000100100: Data = {4'b0101}; //<
    12'b001000100101: Data = {4'b0010}; //+
    12'b001000100110: Data = {4'b0100}; //>
    12'b001000100111: Data = {4'b0100}; //>
    12'b001000101000: Data = {4'b0100}; //>
    12'b001000101001: Data = {4'b0011}; //-
    12'b001000110000: Data = {4'b0111}; //]
    12'b001000110001: Data = {4'b0101}; //<
    12'b001000110010: Data = {4'b0110}; //[
    12'b001000110011: Data = {4'b0100}; //>
    12'b001000110100: Data = {4'b0010}; //+
    12'b001000110101: Data = {4'b0101}; //<
    12'b001000110110: Data = {4'b0011}; //-
    12'b001000110111: Data = {4'b0111}; //]
    12'b001000111000: Data = {4'b0101}; //<
    12'b001000111001: Data = {4'b0010}; //+
    12'b001001000000: Data = {4'b0010}; //+
    12'b001001000001: Data = {4'b0101}; //<
    12'b001001000010: Data = {4'b0101}; //<
    12'b001001000011: Data = {4'b0010}; //+
    12'b001001000100: Data = {4'b0100}; //>
    12'b001001000101: Data = {4'b0100}; //>
    12'b001001000110: Data = {4'b0100}; //>
    12'b001001000111: Data = {4'b0100}; //>
    12'b001001001000: Data = {4'b0100}; //>
    12'b001001001001: Data = {4'b0100}; //>
    12'b001001010000: Data = {4'b0011}; //-
    12'b001001010001: Data = {4'b0111}; //]
    12'b001001010010: Data = {4'b0101}; //<
    12'b001001010011: Data = {4'b0101}; //<
    12'b001001010100: Data = {4'b0110}; //[
    12'b001001010101: Data = {4'b0011}; //-
    12'b001001010110: Data = {4'b0111}; //]
    12'b001001010111: Data = {4'b0101}; //<
    12'b001001011000: Data = {4'b0101}; //<
    12'b001001011001: Data = {4'b0011}; //-
    12'b001001100000: Data = {4'b0101}; //<
    12'b001001100001: Data = {4'b0110}; //[
    12'b001001100010: Data = {4'b0011}; //-
    12'b001001100011: Data = {4'b0100}; //>
    12'b001001100100: Data = {4'b0100}; //>
    12'b001001100101: Data = {4'b0010}; //+
    12'b001001100110: Data = {4'b0101}; //<
    12'b001001100111: Data = {4'b0011}; //-
    12'b001001101000: Data = {4'b0110}; //[
    12'b001001101001: Data = {4'b0100}; //>
    12'b001001110000: Data = {4'b0100}; //>
    12'b001001110001: Data = {4'b0100}; //>
    12'b001001110010: Data = {4'b0111}; //]
    12'b001001110011: Data = {4'b0100}; //>
    12'b001001110100: Data = {4'b0110}; //[
    12'b001001110101: Data = {4'b0110}; //[
    12'b001001110110: Data = {4'b0101}; //<
    12'b001001110111: Data = {4'b0010}; //+
    12'b001001111000: Data = {4'b0100}; //>
    12'b001001111001: Data = {4'b0011}; //-
    12'b001010000000: Data = {4'b0111}; //]
    12'b001010000001: Data = {4'b0100}; //>
    12'b001010000010: Data = {4'b0010}; //+
    12'b001010000011: Data = {4'b0100}; //>
    12'b001010000100: Data = {4'b0100}; //>
    12'b001010000101: Data = {4'b0111}; //]
    12'b001010000110: Data = {4'b0101}; //<
    12'b001010000111: Data = {4'b0101}; //<
    12'b001010001000: Data = {4'b0101}; //<
    12'b001010001001: Data = {4'b0101}; //<
    12'b001010010000: Data = {4'b0101}; //<
    12'b001010010001: Data = {4'b0111}; //]
    12'b001010010010: Data = {4'b0100}; //>
    12'b001010010011: Data = {4'b0110}; //[
    12'b001010010100: Data = {4'b0011}; //-
    12'b001010010101: Data = {4'b0111}; //]
    12'b001010010110: Data = {4'b0100}; //>
    12'b001010010111: Data = {4'b0010}; //+
    12'b001010011000: Data = {4'b0101}; //<
    12'b001010011001: Data = {4'b0101}; //<
    12'b001100000000: Data = {4'b0101}; //<
    12'b001100000001: Data = {4'b0011}; //-
    12'b001100000010: Data = {4'b0110}; //[
    12'b001100000011: Data = {4'b0100}; //>
    12'b001100000100: Data = {4'b0100}; //>
    12'b001100000101: Data = {4'b0010}; //+
    12'b001100000110: Data = {4'b0101}; //<
    12'b001100000111: Data = {4'b0101}; //<
    12'b001100001000: Data = {4'b0011}; //-
    12'b001100001001: Data = {4'b0111}; //]
    12'b001100010000: Data = {4'b0101}; //<
    12'b001100010001: Data = {4'b0111}; //]
    12'b001100010010: Data = {4'b0101}; //<
    12'b001100010011: Data = {4'b0101}; //<
    12'b001100010100: Data = {4'b0101}; //<
    12'b001100010101: Data = {4'b0101}; //<
    12'b001100010110: Data = {4'b0010}; //+
    12'b001100010111: Data = {4'b0100}; //>
    12'b001100011000: Data = {4'b0100}; //>
    12'b001100011001: Data = {4'b0100}; //>
    12'b001100100000: Data = {4'b0100}; //>
    12'b001100100001: Data = {4'b0100}; //>
    12'b001100100010: Data = {4'b0100}; //>
    12'b001100100011: Data = {4'b0100}; //>
    12'b001100100100: Data = {4'b0100}; //>
    12'b001100100101: Data = {4'b0110}; //[
    12'b001100100110: Data = {4'b0011}; //-
    12'b001100100111: Data = {4'b0111}; //]
    12'b001100101000: Data = {4'b0100}; //>
    12'b001100101001: Data = {4'b0110}; //[
    12'b001100110000: Data = {4'b0101}; //<
    12'b001100110001: Data = {4'b0101}; //<
    12'b001100110010: Data = {4'b0101}; //<
    12'b001100110011: Data = {4'b0010}; //+
    12'b001100110100: Data = {4'b0100}; //>
    12'b001100110101: Data = {4'b0100}; //>
    12'b001100110110: Data = {4'b0100}; //>
    12'b001100110111: Data = {4'b0011}; //-
    12'b001100111000: Data = {4'b0111}; //]
    12'b001100111001: Data = {4'b0101}; //<
    12'b001101000000: Data = {4'b0101}; //<
    12'b001101000001: Data = {4'b0010}; //+
    12'b001101000010: Data = {4'b0010}; //+
    12'b001101000011: Data = {4'b0010}; //+
    12'b001101000100: Data = {4'b0010}; //+
    12'b001101000101: Data = {4'b0010}; //+
    12'b001101000110: Data = {4'b0010}; //+
    12'b001101000111: Data = {4'b0010}; //+
    12'b001101001000: Data = {4'b0010}; //+
    12'b001101001001: Data = {4'b0010}; //+
    12'b001101010000: Data = {4'b0010}; //+
    12'b001101010001: Data = {4'b0101}; //<
    12'b001101010010: Data = {4'b0110}; //[
    12'b001101010011: Data = {4'b0011}; //-
    12'b001101010100: Data = {4'b0100}; //>
    12'b001101010101: Data = {4'b0100}; //>
    12'b001101010110: Data = {4'b0010}; //+
    12'b001101010111: Data = {4'b0101}; //<
    12'b001101011000: Data = {4'b0011}; //-
    12'b001101011001: Data = {4'b0110}; //[
    12'b001101100000: Data = {4'b0100}; //>
    12'b001101100001: Data = {4'b0100}; //>
    12'b001101100010: Data = {4'b0100}; //>
    12'b001101100011: Data = {4'b0111}; //]
    12'b001101100100: Data = {4'b0100}; //>
    12'b001101100101: Data = {4'b0110}; //[
    12'b001101100110: Data = {4'b0110}; //[
    12'b001101100111: Data = {4'b0101}; //<
    12'b001101101000: Data = {4'b0010}; //+
    12'b001101101001: Data = {4'b0100}; //>
    12'b001101110000: Data = {4'b0011}; //-
    12'b001101110001: Data = {4'b0111}; //]
    12'b001101110010: Data = {4'b0100}; //>
    12'b001101110011: Data = {4'b0010}; //+
    12'b001101110100: Data = {4'b0100}; //>
    12'b001101110101: Data = {4'b0100}; //>
    12'b001101110110: Data = {4'b0111}; //]
    12'b001101110111: Data = {4'b0101}; //<
    12'b001101111000: Data = {4'b0101}; //<
    12'b001101111001: Data = {4'b0101}; //<
    12'b001110000000: Data = {4'b0101}; //<
    12'b001110000001: Data = {4'b0101}; //<
    12'b001110000010: Data = {4'b0111}; //]
    12'b001110000011: Data = {4'b0100}; //>
    12'b001110000100: Data = {4'b0110}; //[
    12'b001110000101: Data = {4'b0011}; //-
    12'b001110000110: Data = {4'b0111}; //]
    12'b001110000111: Data = {4'b0100}; //>
    12'b001110001000: Data = {4'b0010}; //+
    12'b001110001001: Data = {4'b0100}; //>
    12'b001110010000: Data = {4'b0110}; //[
    12'b001110010001: Data = {4'b0101}; //<
    12'b001110010010: Data = {4'b0101}; //<
    12'b001110010011: Data = {4'b0010}; //+
    12'b001110010100: Data = {4'b0101}; //<
    12'b001110010101: Data = {4'b0010}; //+
    12'b001110010110: Data = {4'b0100}; //>
    12'b001110010111: Data = {4'b0100}; //>
    12'b001110011000: Data = {4'b0100}; //>
    12'b001110011001: Data = {4'b0011}; //-
    12'b010000000000: Data = {4'b0111}; //]
    12'b010000000001: Data = {4'b0101}; //<
    12'b010000000010: Data = {4'b0101}; //<
    12'b010000000011: Data = {4'b0101}; //<
    12'b010000000100: Data = {4'b0101}; //<
    12'b010000000101: Data = {4'b0010}; //+
    12'b010000000110: Data = {4'b0101}; //<
    12'b010000000111: Data = {4'b0010}; //+
    12'b010000001000: Data = {4'b0100}; //>
    12'b010000001001: Data = {4'b0100}; //>
    12'b010000010000: Data = {4'b0110}; //[
    12'b010000010001: Data = {4'b0011}; //-
    12'b010000010010: Data = {4'b0110}; //[
    12'b010000010011: Data = {4'b0011}; //-
    12'b010000010100: Data = {4'b0110}; //[
    12'b010000010101: Data = {4'b0011}; //-
    12'b010000010110: Data = {4'b0110}; //[
    12'b010000010111: Data = {4'b0011}; //-
    12'b010000011000: Data = {4'b0110}; //[
    12'b010000011001: Data = {4'b0011}; //-
    12'b010000100000: Data = {4'b0110}; //[
    12'b010000100001: Data = {4'b0011}; //-
    12'b010000100010: Data = {4'b0110}; //[
    12'b010000100011: Data = {4'b0011}; //-
    12'b010000100100: Data = {4'b0110}; //[
    12'b010000100101: Data = {4'b0011}; //-
    12'b010000100110: Data = {4'b0110}; //[
    12'b010000100111: Data = {4'b0011}; //-
    12'b010000101000: Data = {4'b0101}; //<
    12'b010000101001: Data = {4'b0011}; //-
    12'b010000110000: Data = {4'b0100}; //>
    12'b010000110001: Data = {4'b0110}; //[
    12'b010000110010: Data = {4'b0011}; //-
    12'b010000110011: Data = {4'b0101}; //<
    12'b010000110100: Data = {4'b0010}; //+
    12'b010000110101: Data = {4'b0101}; //<
    12'b010000110110: Data = {4'b0011}; //-
    12'b010000110111: Data = {4'b0100}; //>
    12'b010000111000: Data = {4'b0100}; //>
    12'b010000111001: Data = {4'b0111}; //]
    12'b010001000000: Data = {4'b0111}; //]
    12'b010001000001: Data = {4'b0111}; //]
    12'b010001000010: Data = {4'b0111}; //]
    12'b010001000011: Data = {4'b0111}; //]
    12'b010001000100: Data = {4'b0111}; //]
    12'b010001000101: Data = {4'b0111}; //]
    12'b010001000110: Data = {4'b0111}; //]
    12'b010001000111: Data = {4'b0111}; //]
    12'b010001001000: Data = {4'b0111}; //]
    12'b010001001001: Data = {4'b0101}; //<
    12'b010001010000: Data = {4'b0110}; //[
    12'b010001010001: Data = {4'b0010}; //+
    12'b010001010010: Data = {4'b0010}; //+
    12'b010001010011: Data = {4'b0010}; //+
    12'b010001010100: Data = {4'b0010}; //+
    12'b010001010101: Data = {4'b0010}; //+
    12'b010001010110: Data = {4'b0110}; //[
    12'b010001010111: Data = {4'b0101}; //<
    12'b010001011000: Data = {4'b0101}; //<
    12'b010001011001: Data = {4'b0101}; //<
    12'b010001100000: Data = {4'b0010}; //+
    12'b010001100001: Data = {4'b0010}; //+
    12'b010001100010: Data = {4'b0010}; //+
    12'b010001100011: Data = {4'b0010}; //+
    12'b010001100100: Data = {4'b0010}; //+
    12'b010001100101: Data = {4'b0010}; //+
    12'b010001100110: Data = {4'b0010}; //+
    12'b010001100111: Data = {4'b0010}; //+
    12'b010001101000: Data = {4'b0101}; //<
    12'b010001101001: Data = {4'b0010}; //+
    12'b010001110000: Data = {4'b0010}; //+
    12'b010001110001: Data = {4'b0010}; //+
    12'b010001110010: Data = {4'b0010}; //+
    12'b010001110011: Data = {4'b0010}; //+
    12'b010001110100: Data = {4'b0010}; //+
    12'b010001110101: Data = {4'b0010}; //+
    12'b010001110110: Data = {4'b0010}; //+
    12'b010001110111: Data = {4'b0100}; //>
    12'b010001111000: Data = {4'b0100}; //>
    12'b010001111001: Data = {4'b0100}; //>
    12'b010010000000: Data = {4'b0100}; //>
    12'b010010000001: Data = {4'b0011}; //-
    12'b010010000010: Data = {4'b0111}; //]
    12'b010010000011: Data = {4'b0101}; //<
    12'b010010000100: Data = {4'b0101}; //<
    12'b010010000101: Data = {4'b0101}; //<
    12'b010010000110: Data = {4'b0101}; //<
    12'b010010000111: Data = {4'b0010}; //+
    12'b010010001000: Data = {4'b0101}; //<
    12'b010010001001: Data = {4'b0011}; //-
    12'b010010010000: Data = {4'b0100}; //>
    12'b010010010001: Data = {4'b0100}; //>
    12'b010010010010: Data = {4'b0100}; //>
    12'b010010010011: Data = {4'b0100}; //>
    12'b010010010100: Data = {4'b0110}; //[
    12'b010010010101: Data = {4'b0100}; //>
    12'b010010010110: Data = {4'b0010}; //+
    12'b010010010111: Data = {4'b0101}; //<
    12'b010010011000: Data = {4'b0101}; //<
    12'b010010011001: Data = {4'b0101}; //<
    12'b010100000000: Data = {4'b0010}; //+
    12'b010100000001: Data = {4'b0010}; //+
    12'b010100000010: Data = {4'b0010}; //+
    12'b010100000011: Data = {4'b0010}; //+
    12'b010100000100: Data = {4'b0010}; //+
    12'b010100000101: Data = {4'b0010}; //+
    12'b010100000110: Data = {4'b0010}; //+
    12'b010100000111: Data = {4'b0010}; //+
    12'b010100001000: Data = {4'b0010}; //+
    12'b010100001001: Data = {4'b0101}; //<
    12'b010100010000: Data = {4'b0011}; //-
    12'b010100010001: Data = {4'b0100}; //>
    12'b010100010010: Data = {4'b0100}; //>
    12'b010100010011: Data = {4'b0100}; //>
    12'b010100010100: Data = {4'b0011}; //-
    12'b010100010101: Data = {4'b0111}; //]
    12'b010100010110: Data = {4'b0101}; //<
    12'b010100010111: Data = {4'b0101}; //<
    12'b010100011000: Data = {4'b0101}; //<
    12'b010100011001: Data = {4'b0101}; //<
    12'b010100100000: Data = {4'b0101}; //<
    12'b010100100001: Data = {4'b0110}; //[
    12'b010100100010: Data = {4'b0100}; //>
    12'b010100100011: Data = {4'b0100}; //>
    12'b010100100100: Data = {4'b0010}; //+
    12'b010100100101: Data = {4'b0101}; //<
    12'b010100100110: Data = {4'b0101}; //<
    12'b010100100111: Data = {4'b0011}; //-
    12'b010100101000: Data = {4'b0111}; //]
    12'b010100101001: Data = {4'b0010}; //+
    12'b010100110000: Data = {4'b0101}; //<
    12'b010100110001: Data = {4'b0110}; //[
    12'b010100110010: Data = {4'b0011}; //-
    12'b010100110011: Data = {4'b0100}; //>
    12'b010100110100: Data = {4'b0011}; //-
    12'b010100110101: Data = {4'b0101}; //<
    12'b010100110110: Data = {4'b0111}; //]
    12'b010100110111: Data = {4'b0100}; //>
    12'b010100111000: Data = {4'b0110}; //[
    12'b010100111001: Data = {4'b0100}; //>
    12'b010101000000: Data = {4'b0100}; //>
    12'b010101000001: Data = {4'b1000}; //.
    12'b010101000010: Data = {4'b0101}; //<
    12'b010101000011: Data = {4'b0101}; //<
    12'b010101000100: Data = {4'b0101}; //<
    12'b010101000101: Data = {4'b0101}; //<
    12'b010101000110: Data = {4'b0110}; //[
    12'b010101000111: Data = {4'b0010}; //+
    12'b010101001000: Data = {4'b1000}; //.
    12'b010101001001: Data = {4'b0110}; //[
    12'b010101010000: Data = {4'b0011}; //-
    12'b010101010001: Data = {4'b0111}; //]
    12'b010101010010: Data = {4'b0111}; //]
    12'b010101010011: Data = {4'b0100}; //>
    12'b010101010100: Data = {4'b0100}; //>
    12'b010101010101: Data = {4'b0011}; //-
    12'b010101010110: Data = {4'b0111}; //]
    12'b010101010111: Data = {4'b0100}; //>
    12'b010101011000: Data = {4'b0110}; //[
    12'b010101011001: Data = {4'b0100}; //>
    12'b010101100000: Data = {4'b0100}; //>
    12'b010101100001: Data = {4'b1000}; //.
    12'b010101100010: Data = {4'b0101}; //<
    12'b010101100011: Data = {4'b0101}; //<
    12'b010101100100: Data = {4'b0011}; //-
    12'b010101100101: Data = {4'b0111}; //]
    12'b010101100110: Data = {4'b0100}; //>
    12'b010101100111: Data = {4'b0110}; //[
    12'b010101101000: Data = {4'b0011}; //-
    12'b010101101001: Data = {4'b0111}; //]
    12'b010101110000: Data = {4'b0100}; //>
    12'b010101110001: Data = {4'b0110}; //[
    12'b010101110010: Data = {4'b0011}; //-
    12'b010101110011: Data = {4'b0111}; //]
    12'b010101110100: Data = {4'b0100}; //>
    12'b010101110101: Data = {4'b0100}; //>
    12'b010101110110: Data = {4'b0100}; //>
    12'b010101110111: Data = {4'b0110}; //[
    12'b010101111000: Data = {4'b0100}; //>
    12'b010101111001: Data = {4'b0100}; //>
    12'b010110000000: Data = {4'b0110}; //[
    12'b010110000001: Data = {4'b0101}; //<
    12'b010110000010: Data = {4'b0101}; //<
    12'b010110000011: Data = {4'b0101}; //<
    12'b010110000100: Data = {4'b0101}; //<
    12'b010110000101: Data = {4'b0101}; //<
    12'b010110000110: Data = {4'b0101}; //<
    12'b010110000111: Data = {4'b0101}; //<
    12'b010110001000: Data = {4'b0101}; //<
    12'b010110001001: Data = {4'b0010}; //+
    12'b010110010000: Data = {4'b0100}; //>
    12'b010110010001: Data = {4'b0100}; //>
    12'b010110010010: Data = {4'b0100}; //>
    12'b010110010011: Data = {4'b0100}; //>
    12'b010110010100: Data = {4'b0100}; //>
    12'b010110010101: Data = {4'b0100}; //>
    12'b010110010110: Data = {4'b0100}; //>
    12'b010110010111: Data = {4'b0100}; //>
    12'b010110011000: Data = {4'b0011}; //-
    12'b010110011001: Data = {4'b0111}; //]
    12'b011000000000: Data = {4'b0101}; //<
    12'b011000000001: Data = {4'b0101}; //<
    12'b011000000010: Data = {4'b0011}; //-
    12'b011000000011: Data = {4'b0111}; //]
    12'b011000000100: Data = {4'b0111}; //]
    12'b011000000101: Data = {4'b0100}; //>
    12'b011000000110: Data = {4'b0100}; //>
    12'b011000000111: Data = {4'b0110}; //[
    12'b011000001000: Data = {4'b0011}; //-
    12'b011000001001: Data = {4'b0111}; //]
    12'b011000010000: Data = {4'b0101}; //<
    12'b011000010001: Data = {4'b0101}; //<
    12'b011000010010: Data = {4'b0101}; //<
    12'b011000010011: Data = {4'b0110}; //[
    12'b011000010100: Data = {4'b0011}; //-
    12'b011000010101: Data = {4'b0111}; //]
    12'b011000010110: Data = {4'b0101}; //<
    12'b011000010111: Data = {4'b0101}; //<
    12'b011000011000: Data = {4'b0101}; //<
    12'b011000011001: Data = {4'b0101}; //<
    12'b011000100000: Data = {4'b0101}; //<
    12'b011000100001: Data = {4'b0101}; //<
    12'b011000100010: Data = {4'b0101}; //<
    12'b011000100011: Data = {4'b0101}; //<
    12'b011000100100: Data = {4'b0111}; //]
    12'b011000100101: Data = {4'b0010}; //+
    12'b011000100110: Data = {4'b0010}; //+
    12'b011000100111: Data = {4'b0010}; //+
    12'b011000101000: Data = {4'b0010}; //+
    12'b011000101001: Data = {4'b0010}; //+
    12'b011000110000: Data = {4'b0010}; //+
    12'b011000110001: Data = {4'b0010}; //+
    12'b011000110010: Data = {4'b0010}; //+
    12'b011000110011: Data = {4'b0010}; //+
    12'b011000110100: Data = {4'b0010}; //+
    12'b011000110101: Data = {4'b1000}; //.
    12'b011000110110: Data = {4'b0001}; //H
    12'b011000110111: Data = {4'b0000}; // 
    default: Data = {dataSize{1'bx}};
  endcase

/* verilator lint_on WIDTHEXPAND */
endmodule
