function [7:0] BcdToAscii(
   input [11:0] Bcd
);
  case(Bcd)
    12'h0: BcdToAscii = 8'h0; //  
    12'h1: BcdToAscii = 8'h1; //  
    12'h2: BcdToAscii = 8'h2; //  
    12'h3: BcdToAscii = 8'h3; //  
    12'h4: BcdToAscii = 8'h4; //  
    12'h5: BcdToAscii = 8'h5; //  
    12'h6: BcdToAscii = 8'h6; //  
    12'h7: BcdToAscii = 8'h7; //  
    12'h8: BcdToAscii = 8'h8; //  
    12'h9: BcdToAscii = 8'h9; //  
    12'h10: BcdToAscii = 8'ha; //  
    12'h11: BcdToAscii = 8'hb; //  
    12'h12: BcdToAscii = 8'hc; //  
    12'h13: BcdToAscii = 8'hd; //  
    12'h14: BcdToAscii = 8'he; //  
    12'h15: BcdToAscii = 8'hf; //  
    12'h16: BcdToAscii = 8'h10; //  
    12'h17: BcdToAscii = 8'h11; //  
    12'h18: BcdToAscii = 8'h12; //  
    12'h19: BcdToAscii = 8'h13; //  
    12'h20: BcdToAscii = 8'h14; //  
    12'h21: BcdToAscii = 8'h15; //  
    12'h22: BcdToAscii = 8'h16; //  
    12'h23: BcdToAscii = 8'h17; //  
    12'h24: BcdToAscii = 8'h18; //  
    12'h25: BcdToAscii = 8'h19; //  
    12'h26: BcdToAscii = 8'h1a; //  
    12'h27: BcdToAscii = 8'h1b; //  
    12'h28: BcdToAscii = 8'h1c; //  
    12'h29: BcdToAscii = 8'h1d; //  
    12'h30: BcdToAscii = 8'h1e; //  
    12'h31: BcdToAscii = 8'h1f; //  
    12'h32: BcdToAscii = 8'h20; //  
    12'h33: BcdToAscii = 8'h21; //! 
    12'h34: BcdToAscii = 8'h22; //" 
    12'h35: BcdToAscii = 8'h23; //# 
    12'h36: BcdToAscii = 8'h24; //$ 
    12'h37: BcdToAscii = 8'h25; //% 
    12'h38: BcdToAscii = 8'h26; //& 
    12'h39: BcdToAscii = 8'h27; //' 
    12'h40: BcdToAscii = 8'h28; //( 
    12'h41: BcdToAscii = 8'h29; //) 
    12'h42: BcdToAscii = 8'h2a; //* 
    12'h43: BcdToAscii = 8'h2b; //+ 
    12'h44: BcdToAscii = 8'h2c; //, 
    12'h45: BcdToAscii = 8'h2d; //- 
    12'h46: BcdToAscii = 8'h2e; //. 
    12'h47: BcdToAscii = 8'h2f; /// 
    12'h48: BcdToAscii = 8'h30; //0 
    12'h49: BcdToAscii = 8'h31; //1 
    12'h50: BcdToAscii = 8'h32; //2 
    12'h51: BcdToAscii = 8'h33; //3 
    12'h52: BcdToAscii = 8'h34; //4 
    12'h53: BcdToAscii = 8'h35; //5 
    12'h54: BcdToAscii = 8'h36; //6 
    12'h55: BcdToAscii = 8'h37; //7 
    12'h56: BcdToAscii = 8'h38; //8 
    12'h57: BcdToAscii = 8'h39; //9 
    12'h58: BcdToAscii = 8'h3a; //: 
    12'h59: BcdToAscii = 8'h3b; //; 
    12'h60: BcdToAscii = 8'h3c; //< 
    12'h61: BcdToAscii = 8'h3d; //= 
    12'h62: BcdToAscii = 8'h3e; //> 
    12'h63: BcdToAscii = 8'h3f; //? 
    12'h64: BcdToAscii = 8'h40; //@ 
    12'h65: BcdToAscii = 8'h41; //A 
    12'h66: BcdToAscii = 8'h42; //B 
    12'h67: BcdToAscii = 8'h43; //C 
    12'h68: BcdToAscii = 8'h44; //D 
    12'h69: BcdToAscii = 8'h45; //E 
    12'h70: BcdToAscii = 8'h46; //F 
    12'h71: BcdToAscii = 8'h47; //G 
    12'h72: BcdToAscii = 8'h48; //H 
    12'h73: BcdToAscii = 8'h49; //I 
    12'h74: BcdToAscii = 8'h4a; //J 
    12'h75: BcdToAscii = 8'h4b; //K 
    12'h76: BcdToAscii = 8'h4c; //L 
    12'h77: BcdToAscii = 8'h4d; //M 
    12'h78: BcdToAscii = 8'h4e; //N 
    12'h79: BcdToAscii = 8'h4f; //O 
    12'h80: BcdToAscii = 8'h50; //P 
    12'h81: BcdToAscii = 8'h51; //Q 
    12'h82: BcdToAscii = 8'h52; //R 
    12'h83: BcdToAscii = 8'h53; //S 
    12'h84: BcdToAscii = 8'h54; //T 
    12'h85: BcdToAscii = 8'h55; //U 
    12'h86: BcdToAscii = 8'h56; //V 
    12'h87: BcdToAscii = 8'h57; //W 
    12'h88: BcdToAscii = 8'h58; //X 
    12'h89: BcdToAscii = 8'h59; //Y 
    12'h90: BcdToAscii = 8'h5a; //Z 
    12'h91: BcdToAscii = 8'h5b; //[ 
    12'h92: BcdToAscii = 8'h5c; //\ 
    12'h93: BcdToAscii = 8'h5d; //] 
    12'h94: BcdToAscii = 8'h5e; //^ 
    12'h95: BcdToAscii = 8'h5f; //_ 
    12'h96: BcdToAscii = 8'h60; //` 
    12'h97: BcdToAscii = 8'h61; //a 
    12'h98: BcdToAscii = 8'h62; //b 
    12'h99: BcdToAscii = 8'h63; //c 
    12'h100: BcdToAscii = 8'h64; //d 
    12'h101: BcdToAscii = 8'h65; //e 
    12'h102: BcdToAscii = 8'h66; //f 
    12'h103: BcdToAscii = 8'h67; //g 
    12'h104: BcdToAscii = 8'h68; //h 
    12'h105: BcdToAscii = 8'h69; //i 
    12'h106: BcdToAscii = 8'h6a; //j 
    12'h107: BcdToAscii = 8'h6b; //k 
    12'h108: BcdToAscii = 8'h6c; //l 
    12'h109: BcdToAscii = 8'h6d; //m 
    12'h110: BcdToAscii = 8'h6e; //n 
    12'h111: BcdToAscii = 8'h6f; //o 
    12'h112: BcdToAscii = 8'h70; //p 
    12'h113: BcdToAscii = 8'h71; //q 
    12'h114: BcdToAscii = 8'h72; //r 
    12'h115: BcdToAscii = 8'h73; //s 
    12'h116: BcdToAscii = 8'h74; //t 
    12'h117: BcdToAscii = 8'h75; //u 
    12'h118: BcdToAscii = 8'h76; //v 
    12'h119: BcdToAscii = 8'h77; //w 
    12'h120: BcdToAscii = 8'h78; //x 
    12'h121: BcdToAscii = 8'h79; //y 
    12'h122: BcdToAscii = 8'h7a; //z 
    12'h123: BcdToAscii = 8'h7b; //{ 
    12'h124: BcdToAscii = 8'h7c; //| 
    12'h125: BcdToAscii = 8'h7d; //} 
    12'h126: BcdToAscii = 8'h7e; //~ 
    12'h127: BcdToAscii = 8'h7f; // 
    12'h128: BcdToAscii = 8'h80; // 
    12'h129: BcdToAscii = 8'h81; // 
    12'h130: BcdToAscii = 8'h82; // 
    12'h131: BcdToAscii = 8'h83; // 
    12'h132: BcdToAscii = 8'h84; // 
    12'h133: BcdToAscii = 8'h85; // 
    12'h134: BcdToAscii = 8'h86; // 
    12'h135: BcdToAscii = 8'h87; // 
    12'h136: BcdToAscii = 8'h88; // 
    12'h137: BcdToAscii = 8'h89; // 
    12'h138: BcdToAscii = 8'h8a; // 
    12'h139: BcdToAscii = 8'h8b; // 
    12'h140: BcdToAscii = 8'h8c; // 
    12'h141: BcdToAscii = 8'h8d; // 
    12'h142: BcdToAscii = 8'h8e; // 
    12'h143: BcdToAscii = 8'h8f; // 
    12'h144: BcdToAscii = 8'h90; // 
    12'h145: BcdToAscii = 8'h91; // 
    12'h146: BcdToAscii = 8'h92; // 
    12'h147: BcdToAscii = 8'h93; // 
    12'h148: BcdToAscii = 8'h94; // 
    12'h149: BcdToAscii = 8'h95; // 
    12'h150: BcdToAscii = 8'h96; // 
    12'h151: BcdToAscii = 8'h97; // 
    12'h152: BcdToAscii = 8'h98; // 
    12'h153: BcdToAscii = 8'h99; // 
    12'h154: BcdToAscii = 8'h9a; // 
    12'h155: BcdToAscii = 8'h9b; // 
    12'h156: BcdToAscii = 8'h9c; // 
    12'h157: BcdToAscii = 8'h9d; // 
    12'h158: BcdToAscii = 8'h9e; // 
    12'h159: BcdToAscii = 8'h9f; // 
    12'h160: BcdToAscii = 8'ha0; //  
    12'h161: BcdToAscii = 8'ha1; //¡ 
    12'h162: BcdToAscii = 8'ha2; //¢ 
    12'h163: BcdToAscii = 8'ha3; //£ 
    12'h164: BcdToAscii = 8'ha4; //¤ 
    12'h165: BcdToAscii = 8'ha5; //¥ 
    12'h166: BcdToAscii = 8'ha6; //¦ 
    12'h167: BcdToAscii = 8'ha7; //§ 
    12'h168: BcdToAscii = 8'ha8; //¨ 
    12'h169: BcdToAscii = 8'ha9; //© 
    12'h170: BcdToAscii = 8'haa; //ª 
    12'h171: BcdToAscii = 8'hab; //« 
    12'h172: BcdToAscii = 8'hac; //¬ 
    12'h173: BcdToAscii = 8'had; //­ 
    12'h174: BcdToAscii = 8'hae; //® 
    12'h175: BcdToAscii = 8'haf; //¯ 
    12'h176: BcdToAscii = 8'hb0; //° 
    12'h177: BcdToAscii = 8'hb1; //± 
    12'h178: BcdToAscii = 8'hb2; //² 
    12'h179: BcdToAscii = 8'hb3; //³ 
    12'h180: BcdToAscii = 8'hb4; //´ 
    12'h181: BcdToAscii = 8'hb5; //µ 
    12'h182: BcdToAscii = 8'hb6; //¶ 
    12'h183: BcdToAscii = 8'hb7; //· 
    12'h184: BcdToAscii = 8'hb8; //¸ 
    12'h185: BcdToAscii = 8'hb9; //¹ 
    12'h186: BcdToAscii = 8'hba; //º 
    12'h187: BcdToAscii = 8'hbb; //» 
    12'h188: BcdToAscii = 8'hbc; //¼ 
    12'h189: BcdToAscii = 8'hbd; //½ 
    12'h190: BcdToAscii = 8'hbe; //¾ 
    12'h191: BcdToAscii = 8'hbf; //¿ 
    12'h192: BcdToAscii = 8'hc0; //À 
    12'h193: BcdToAscii = 8'hc1; //Á 
    12'h194: BcdToAscii = 8'hc2; //Â 
    12'h195: BcdToAscii = 8'hc3; //Ã 
    12'h196: BcdToAscii = 8'hc4; //Ä 
    12'h197: BcdToAscii = 8'hc5; //Å 
    12'h198: BcdToAscii = 8'hc6; //Æ 
    12'h199: BcdToAscii = 8'hc7; //Ç 
    12'h200: BcdToAscii = 8'hc8; //È 
    12'h201: BcdToAscii = 8'hc9; //É 
    12'h202: BcdToAscii = 8'hca; //Ê 
    12'h203: BcdToAscii = 8'hcb; //Ë 
    12'h204: BcdToAscii = 8'hcc; //Ì 
    12'h205: BcdToAscii = 8'hcd; //Í 
    12'h206: BcdToAscii = 8'hce; //Î 
    12'h207: BcdToAscii = 8'hcf; //Ï 
    12'h208: BcdToAscii = 8'hd0; //Ð 
    12'h209: BcdToAscii = 8'hd1; //Ñ 
    12'h210: BcdToAscii = 8'hd2; //Ò 
    12'h211: BcdToAscii = 8'hd3; //Ó 
    12'h212: BcdToAscii = 8'hd4; //Ô 
    12'h213: BcdToAscii = 8'hd5; //Õ 
    12'h214: BcdToAscii = 8'hd6; //Ö 
    12'h215: BcdToAscii = 8'hd7; //× 
    12'h216: BcdToAscii = 8'hd8; //Ø 
    12'h217: BcdToAscii = 8'hd9; //Ù 
    12'h218: BcdToAscii = 8'hda; //Ú 
    12'h219: BcdToAscii = 8'hdb; //Û 
    12'h220: BcdToAscii = 8'hdc; //Ü 
    12'h221: BcdToAscii = 8'hdd; //Ý 
    12'h222: BcdToAscii = 8'hde; //Þ 
    12'h223: BcdToAscii = 8'hdf; //ß 
    12'h224: BcdToAscii = 8'he0; //à 
    12'h225: BcdToAscii = 8'he1; //á 
    12'h226: BcdToAscii = 8'he2; //â 
    12'h227: BcdToAscii = 8'he3; //ã 
    12'h228: BcdToAscii = 8'he4; //ä 
    12'h229: BcdToAscii = 8'he5; //å 
    12'h230: BcdToAscii = 8'he6; //æ 
    12'h231: BcdToAscii = 8'he7; //ç 
    12'h232: BcdToAscii = 8'he8; //è 
    12'h233: BcdToAscii = 8'he9; //é 
    12'h234: BcdToAscii = 8'hea; //ê 
    12'h235: BcdToAscii = 8'heb; //ë 
    12'h236: BcdToAscii = 8'hec; //ì 
    12'h237: BcdToAscii = 8'hed; //í 
    12'h238: BcdToAscii = 8'hee; //î 
    12'h239: BcdToAscii = 8'hef; //ï 
    12'h240: BcdToAscii = 8'hf0; //ð 
    12'h241: BcdToAscii = 8'hf1; //ñ 
    12'h242: BcdToAscii = 8'hf2; //ò 
    12'h243: BcdToAscii = 8'hf3; //ó 
    12'h244: BcdToAscii = 8'hf4; //ô 
    12'h245: BcdToAscii = 8'hf5; //õ 
    12'h246: BcdToAscii = 8'hf6; //ö 
    12'h247: BcdToAscii = 8'hf7; //÷ 
    12'h248: BcdToAscii = 8'hf8; //ø 
    12'h249: BcdToAscii = 8'hf9; //ù 
    12'h250: BcdToAscii = 8'hfa; //ú 
    12'h251: BcdToAscii = 8'hfb; //û 
    12'h252: BcdToAscii = 8'hfc; //ü 
    12'h253: BcdToAscii = 8'hfd; //ý 
    12'h254: BcdToAscii = 8'hfe; //þ 
    12'h255: BcdToAscii = 8'hff; //ÿ 
    default: BcdToAscii = {8'bx};
  endcase
endfunction
