module IpBlock();


endmodule;