function [11:0] AsciiToBcd(
   input [7:0] ascii
);
  case(ascii)
    8'h0: AsciiToBcd = 12'h0; //  
    8'h1: AsciiToBcd = 12'h1; //  
    8'h2: AsciiToBcd = 12'h2; //  
    8'h3: AsciiToBcd = 12'h3; //  
    8'h4: AsciiToBcd = 12'h4; //  
    8'h5: AsciiToBcd = 12'h5; //  
    8'h6: AsciiToBcd = 12'h6; //  
    8'h7: AsciiToBcd = 12'h7; //  
    8'h8: AsciiToBcd = 12'h8; //  
    8'h9: AsciiToBcd = 12'h9; //  
    8'h10: AsciiToBcd = 12'ha; //  
    8'h11: AsciiToBcd = 12'hb; //  
    8'h12: AsciiToBcd = 12'hc; //  
    8'h13: AsciiToBcd = 12'hd; //  
    8'h14: AsciiToBcd = 12'he; //  
    8'h15: AsciiToBcd = 12'hf; //  
    8'h16: AsciiToBcd = 12'h10; //  
    8'h17: AsciiToBcd = 12'h11; //  
    8'h18: AsciiToBcd = 12'h12; //  
    8'h19: AsciiToBcd = 12'h13; //  
    8'h20: AsciiToBcd = 12'h14; //  
    8'h21: AsciiToBcd = 12'h15; //  
    8'h22: AsciiToBcd = 12'h16; //  
    8'h23: AsciiToBcd = 12'h17; //  
    8'h24: AsciiToBcd = 12'h18; //  
    8'h25: AsciiToBcd = 12'h19; //  
    8'h26: AsciiToBcd = 12'h1a; //  
    8'h27: AsciiToBcd = 12'h1b; //  
    8'h28: AsciiToBcd = 12'h1c; //  
    8'h29: AsciiToBcd = 12'h1d; //  
    8'h30: AsciiToBcd = 12'h1e; //  
    8'h31: AsciiToBcd = 12'h1f; //  
    8'h32: AsciiToBcd = 12'h20; //  
    8'h33: AsciiToBcd = 12'h21; //! 
    8'h34: AsciiToBcd = 12'h22; //" 
    8'h35: AsciiToBcd = 12'h23; //# 
    8'h36: AsciiToBcd = 12'h24; //$ 
    8'h37: AsciiToBcd = 12'h25; //% 
    8'h38: AsciiToBcd = 12'h26; //& 
    8'h39: AsciiToBcd = 12'h27; //' 
    8'h40: AsciiToBcd = 12'h28; //( 
    8'h41: AsciiToBcd = 12'h29; //) 
    8'h42: AsciiToBcd = 12'h2a; //* 
    8'h43: AsciiToBcd = 12'h2b; //+ 
    8'h44: AsciiToBcd = 12'h2c; //, 
    8'h45: AsciiToBcd = 12'h2d; //- 
    8'h46: AsciiToBcd = 12'h2e; //. 
    8'h47: AsciiToBcd = 12'h2f; /// 
    8'h48: AsciiToBcd = 12'h30; //0 
    8'h49: AsciiToBcd = 12'h31; //1 
    8'h50: AsciiToBcd = 12'h32; //2 
    8'h51: AsciiToBcd = 12'h33; //3 
    8'h52: AsciiToBcd = 12'h34; //4 
    8'h53: AsciiToBcd = 12'h35; //5 
    8'h54: AsciiToBcd = 12'h36; //6 
    8'h55: AsciiToBcd = 12'h37; //7 
    8'h56: AsciiToBcd = 12'h38; //8 
    8'h57: AsciiToBcd = 12'h39; //9 
    8'h58: AsciiToBcd = 12'h3a; //: 
    8'h59: AsciiToBcd = 12'h3b; //; 
    8'h60: AsciiToBcd = 12'h3c; //< 
    8'h61: AsciiToBcd = 12'h3d; //= 
    8'h62: AsciiToBcd = 12'h3e; //> 
    8'h63: AsciiToBcd = 12'h3f; //? 
    8'h64: AsciiToBcd = 12'h40; //@ 
    8'h65: AsciiToBcd = 12'h41; //A 
    8'h66: AsciiToBcd = 12'h42; //B 
    8'h67: AsciiToBcd = 12'h43; //C 
    8'h68: AsciiToBcd = 12'h44; //D 
    8'h69: AsciiToBcd = 12'h45; //E 
    8'h70: AsciiToBcd = 12'h46; //F 
    8'h71: AsciiToBcd = 12'h47; //G 
    8'h72: AsciiToBcd = 12'h48; //H 
    8'h73: AsciiToBcd = 12'h49; //I 
    8'h74: AsciiToBcd = 12'h4a; //J 
    8'h75: AsciiToBcd = 12'h4b; //K 
    8'h76: AsciiToBcd = 12'h4c; //L 
    8'h77: AsciiToBcd = 12'h4d; //M 
    8'h78: AsciiToBcd = 12'h4e; //N 
    8'h79: AsciiToBcd = 12'h4f; //O 
    8'h80: AsciiToBcd = 12'h50; //P 
    8'h81: AsciiToBcd = 12'h51; //Q 
    8'h82: AsciiToBcd = 12'h52; //R 
    8'h83: AsciiToBcd = 12'h53; //S 
    8'h84: AsciiToBcd = 12'h54; //T 
    8'h85: AsciiToBcd = 12'h55; //U 
    8'h86: AsciiToBcd = 12'h56; //V 
    8'h87: AsciiToBcd = 12'h57; //W 
    8'h88: AsciiToBcd = 12'h58; //X 
    8'h89: AsciiToBcd = 12'h59; //Y 
    8'h90: AsciiToBcd = 12'h5a; //Z 
    8'h91: AsciiToBcd = 12'h5b; //[ 
    8'h92: AsciiToBcd = 12'h5c; //\ 
    8'h93: AsciiToBcd = 12'h5d; //] 
    8'h94: AsciiToBcd = 12'h5e; //^ 
    8'h95: AsciiToBcd = 12'h5f; //_ 
    8'h96: AsciiToBcd = 12'h60; //` 
    8'h97: AsciiToBcd = 12'h61; //a 
    8'h98: AsciiToBcd = 12'h62; //b 
    8'h99: AsciiToBcd = 12'h63; //c 
    8'h100: AsciiToBcd = 12'h64; //d 
    8'h101: AsciiToBcd = 12'h65; //e 
    8'h102: AsciiToBcd = 12'h66; //f 
    8'h103: AsciiToBcd = 12'h67; //g 
    8'h104: AsciiToBcd = 12'h68; //h 
    8'h105: AsciiToBcd = 12'h69; //i 
    8'h106: AsciiToBcd = 12'h6a; //j 
    8'h107: AsciiToBcd = 12'h6b; //k 
    8'h108: AsciiToBcd = 12'h6c; //l 
    8'h109: AsciiToBcd = 12'h6d; //m 
    8'h110: AsciiToBcd = 12'h6e; //n 
    8'h111: AsciiToBcd = 12'h6f; //o 
    8'h112: AsciiToBcd = 12'h70; //p 
    8'h113: AsciiToBcd = 12'h71; //q 
    8'h114: AsciiToBcd = 12'h72; //r 
    8'h115: AsciiToBcd = 12'h73; //s 
    8'h116: AsciiToBcd = 12'h74; //t 
    8'h117: AsciiToBcd = 12'h75; //u 
    8'h118: AsciiToBcd = 12'h76; //v 
    8'h119: AsciiToBcd = 12'h77; //w 
    8'h120: AsciiToBcd = 12'h78; //x 
    8'h121: AsciiToBcd = 12'h79; //y 
    8'h122: AsciiToBcd = 12'h7a; //z 
    8'h123: AsciiToBcd = 12'h7b; //{ 
    8'h124: AsciiToBcd = 12'h7c; //| 
    8'h125: AsciiToBcd = 12'h7d; //} 
    8'h126: AsciiToBcd = 12'h7e; //~ 
    8'h127: AsciiToBcd = 12'h7f; // 
    8'h128: AsciiToBcd = 12'h80; // 
    8'h129: AsciiToBcd = 12'h81; // 
    8'h130: AsciiToBcd = 12'h82; // 
    8'h131: AsciiToBcd = 12'h83; // 
    8'h132: AsciiToBcd = 12'h84; // 
    8'h133: AsciiToBcd = 12'h85; // 
    8'h134: AsciiToBcd = 12'h86; // 
    8'h135: AsciiToBcd = 12'h87; // 
    8'h136: AsciiToBcd = 12'h88; // 
    8'h137: AsciiToBcd = 12'h89; // 
    8'h138: AsciiToBcd = 12'h8a; // 
    8'h139: AsciiToBcd = 12'h8b; // 
    8'h140: AsciiToBcd = 12'h8c; // 
    8'h141: AsciiToBcd = 12'h8d; // 
    8'h142: AsciiToBcd = 12'h8e; // 
    8'h143: AsciiToBcd = 12'h8f; // 
    8'h144: AsciiToBcd = 12'h90; // 
    8'h145: AsciiToBcd = 12'h91; // 
    8'h146: AsciiToBcd = 12'h92; // 
    8'h147: AsciiToBcd = 12'h93; // 
    8'h148: AsciiToBcd = 12'h94; // 
    8'h149: AsciiToBcd = 12'h95; // 
    8'h150: AsciiToBcd = 12'h96; // 
    8'h151: AsciiToBcd = 12'h97; // 
    8'h152: AsciiToBcd = 12'h98; // 
    8'h153: AsciiToBcd = 12'h99; // 
    8'h154: AsciiToBcd = 12'h9a; // 
    8'h155: AsciiToBcd = 12'h9b; // 
    8'h156: AsciiToBcd = 12'h9c; // 
    8'h157: AsciiToBcd = 12'h9d; // 
    8'h158: AsciiToBcd = 12'h9e; // 
    8'h159: AsciiToBcd = 12'h9f; // 
    8'h160: AsciiToBcd = 12'ha0; //  
    8'h161: AsciiToBcd = 12'ha1; //¡ 
    8'h162: AsciiToBcd = 12'ha2; //¢ 
    8'h163: AsciiToBcd = 12'ha3; //£ 
    8'h164: AsciiToBcd = 12'ha4; //¤ 
    8'h165: AsciiToBcd = 12'ha5; //¥ 
    8'h166: AsciiToBcd = 12'ha6; //¦ 
    8'h167: AsciiToBcd = 12'ha7; //§ 
    8'h168: AsciiToBcd = 12'ha8; //¨ 
    8'h169: AsciiToBcd = 12'ha9; //© 
    8'h170: AsciiToBcd = 12'haa; //ª 
    8'h171: AsciiToBcd = 12'hab; //« 
    8'h172: AsciiToBcd = 12'hac; //¬ 
    8'h173: AsciiToBcd = 12'had; //­ 
    8'h174: AsciiToBcd = 12'hae; //® 
    8'h175: AsciiToBcd = 12'haf; //¯ 
    8'h176: AsciiToBcd = 12'hb0; //° 
    8'h177: AsciiToBcd = 12'hb1; //± 
    8'h178: AsciiToBcd = 12'hb2; //² 
    8'h179: AsciiToBcd = 12'hb3; //³ 
    8'h180: AsciiToBcd = 12'hb4; //´ 
    8'h181: AsciiToBcd = 12'hb5; //µ 
    8'h182: AsciiToBcd = 12'hb6; //¶ 
    8'h183: AsciiToBcd = 12'hb7; //· 
    8'h184: AsciiToBcd = 12'hb8; //¸ 
    8'h185: AsciiToBcd = 12'hb9; //¹ 
    8'h186: AsciiToBcd = 12'hba; //º 
    8'h187: AsciiToBcd = 12'hbb; //» 
    8'h188: AsciiToBcd = 12'hbc; //¼ 
    8'h189: AsciiToBcd = 12'hbd; //½ 
    8'h190: AsciiToBcd = 12'hbe; //¾ 
    8'h191: AsciiToBcd = 12'hbf; //¿ 
    8'h192: AsciiToBcd = 12'hc0; //À 
    8'h193: AsciiToBcd = 12'hc1; //Á 
    8'h194: AsciiToBcd = 12'hc2; //Â 
    8'h195: AsciiToBcd = 12'hc3; //Ã 
    8'h196: AsciiToBcd = 12'hc4; //Ä 
    8'h197: AsciiToBcd = 12'hc5; //Å 
    8'h198: AsciiToBcd = 12'hc6; //Æ 
    8'h199: AsciiToBcd = 12'hc7; //Ç 
    8'h200: AsciiToBcd = 12'hc8; //È 
    8'h201: AsciiToBcd = 12'hc9; //É 
    8'h202: AsciiToBcd = 12'hca; //Ê 
    8'h203: AsciiToBcd = 12'hcb; //Ë 
    8'h204: AsciiToBcd = 12'hcc; //Ì 
    8'h205: AsciiToBcd = 12'hcd; //Í 
    8'h206: AsciiToBcd = 12'hce; //Î 
    8'h207: AsciiToBcd = 12'hcf; //Ï 
    8'h208: AsciiToBcd = 12'hd0; //Ð 
    8'h209: AsciiToBcd = 12'hd1; //Ñ 
    8'h210: AsciiToBcd = 12'hd2; //Ò 
    8'h211: AsciiToBcd = 12'hd3; //Ó 
    8'h212: AsciiToBcd = 12'hd4; //Ô 
    8'h213: AsciiToBcd = 12'hd5; //Õ 
    8'h214: AsciiToBcd = 12'hd6; //Ö 
    8'h215: AsciiToBcd = 12'hd7; //× 
    8'h216: AsciiToBcd = 12'hd8; //Ø 
    8'h217: AsciiToBcd = 12'hd9; //Ù 
    8'h218: AsciiToBcd = 12'hda; //Ú 
    8'h219: AsciiToBcd = 12'hdb; //Û 
    8'h220: AsciiToBcd = 12'hdc; //Ü 
    8'h221: AsciiToBcd = 12'hdd; //Ý 
    8'h222: AsciiToBcd = 12'hde; //Þ 
    8'h223: AsciiToBcd = 12'hdf; //ß 
    8'h224: AsciiToBcd = 12'he0; //à 
    8'h225: AsciiToBcd = 12'he1; //á 
    8'h226: AsciiToBcd = 12'he2; //â 
    8'h227: AsciiToBcd = 12'he3; //ã 
    8'h228: AsciiToBcd = 12'he4; //ä 
    8'h229: AsciiToBcd = 12'he5; //å 
    8'h230: AsciiToBcd = 12'he6; //æ 
    8'h231: AsciiToBcd = 12'he7; //ç 
    8'h232: AsciiToBcd = 12'he8; //è 
    8'h233: AsciiToBcd = 12'he9; //é 
    8'h234: AsciiToBcd = 12'hea; //ê 
    8'h235: AsciiToBcd = 12'heb; //ë 
    8'h236: AsciiToBcd = 12'hec; //ì 
    8'h237: AsciiToBcd = 12'hed; //í 
    8'h238: AsciiToBcd = 12'hee; //î 
    8'h239: AsciiToBcd = 12'hef; //ï 
    8'h240: AsciiToBcd = 12'hf0; //ð 
    8'h241: AsciiToBcd = 12'hf1; //ñ 
    8'h242: AsciiToBcd = 12'hf2; //ò 
    8'h243: AsciiToBcd = 12'hf3; //ó 
    8'h244: AsciiToBcd = 12'hf4; //ô 
    8'h245: AsciiToBcd = 12'hf5; //õ 
    8'h246: AsciiToBcd = 12'hf6; //ö 
    8'h247: AsciiToBcd = 12'hf7; //÷ 
    8'h248: AsciiToBcd = 12'hf8; //ø 
    8'h249: AsciiToBcd = 12'hf9; //ù 
    8'h250: AsciiToBcd = 12'hfa; //ú 
    8'h251: AsciiToBcd = 12'hfb; //û 
    8'h252: AsciiToBcd = 12'hfc; //ü 
    8'h253: AsciiToBcd = 12'hfd; //ý 
    8'h254: AsciiToBcd = 12'hfe; //þ 
    8'h255: AsciiToBcd = 12'hff; //ÿ 
    default: AsciiToBcd = {12'bx};n  endcase
endfunction
