function [7:0] BcdToAscii(
   input [12:0] Bcd
);
  case(Bdc)
    12'h0: BcdToAscii = 8'h0; //  
    12'h1: BcdToAscii = 8'h1; //  
    12'h2: BcdToAscii = 8'h2; //  
    12'h3: BcdToAscii = 8'h3; //  
    12'h4: BcdToAscii = 8'h4; //  
    12'h5: BcdToAscii = 8'h5; //  
    12'h6: BcdToAscii = 8'h6; //  
    12'h7: BcdToAscii = 8'h7; //  
    12'h8: BcdToAscii = 8'h8; //  
    12'h9: BcdToAscii = 8'h9; //  
    12'ha: BcdToAscii = 8'h10; //  
    12'hb: BcdToAscii = 8'h11; //  
    12'hc: BcdToAscii = 8'h12; //  
    12'hd: BcdToAscii = 8'h13; //  
    12'he: BcdToAscii = 8'h14; //  
    12'hf: BcdToAscii = 8'h15; //  
    12'h10: BcdToAscii = 8'h16; //  
    12'h11: BcdToAscii = 8'h17; //  
    12'h12: BcdToAscii = 8'h18; //  
    12'h13: BcdToAscii = 8'h19; //  
    12'h14: BcdToAscii = 8'h20; //  
    12'h15: BcdToAscii = 8'h21; //  
    12'h16: BcdToAscii = 8'h22; //  
    12'h17: BcdToAscii = 8'h23; //  
    12'h18: BcdToAscii = 8'h24; //  
    12'h19: BcdToAscii = 8'h25; //  
    12'h1a: BcdToAscii = 8'h26; //  
    12'h1b: BcdToAscii = 8'h27; //  
    12'h1c: BcdToAscii = 8'h28; //  
    12'h1d: BcdToAscii = 8'h29; //  
    12'h1e: BcdToAscii = 8'h30; //  
    12'h1f: BcdToAscii = 8'h31; //  
    12'h20: BcdToAscii = 8'h32; //  
    12'h21: BcdToAscii = 8'h33; //! 
    12'h22: BcdToAscii = 8'h34; //" 
    12'h23: BcdToAscii = 8'h35; //# 
    12'h24: BcdToAscii = 8'h36; //$ 
    12'h25: BcdToAscii = 8'h37; //% 
    12'h26: BcdToAscii = 8'h38; //& 
    12'h27: BcdToAscii = 8'h39; //' 
    12'h28: BcdToAscii = 8'h40; //( 
    12'h29: BcdToAscii = 8'h41; //) 
    12'h2a: BcdToAscii = 8'h42; //* 
    12'h2b: BcdToAscii = 8'h43; //+ 
    12'h2c: BcdToAscii = 8'h44; //, 
    12'h2d: BcdToAscii = 8'h45; //- 
    12'h2e: BcdToAscii = 8'h46; //. 
    12'h2f: BcdToAscii = 8'h47; /// 
    12'h30: BcdToAscii = 8'h48; //0 
    12'h31: BcdToAscii = 8'h49; //1 
    12'h32: BcdToAscii = 8'h50; //2 
    12'h33: BcdToAscii = 8'h51; //3 
    12'h34: BcdToAscii = 8'h52; //4 
    12'h35: BcdToAscii = 8'h53; //5 
    12'h36: BcdToAscii = 8'h54; //6 
    12'h37: BcdToAscii = 8'h55; //7 
    12'h38: BcdToAscii = 8'h56; //8 
    12'h39: BcdToAscii = 8'h57; //9 
    12'h3a: BcdToAscii = 8'h58; //: 
    12'h3b: BcdToAscii = 8'h59; //; 
    12'h3c: BcdToAscii = 8'h60; //< 
    12'h3d: BcdToAscii = 8'h61; //= 
    12'h3e: BcdToAscii = 8'h62; //> 
    12'h3f: BcdToAscii = 8'h63; //? 
    12'h40: BcdToAscii = 8'h64; //@ 
    12'h41: BcdToAscii = 8'h65; //A 
    12'h42: BcdToAscii = 8'h66; //B 
    12'h43: BcdToAscii = 8'h67; //C 
    12'h44: BcdToAscii = 8'h68; //D 
    12'h45: BcdToAscii = 8'h69; //E 
    12'h46: BcdToAscii = 8'h70; //F 
    12'h47: BcdToAscii = 8'h71; //G 
    12'h48: BcdToAscii = 8'h72; //H 
    12'h49: BcdToAscii = 8'h73; //I 
    12'h4a: BcdToAscii = 8'h74; //J 
    12'h4b: BcdToAscii = 8'h75; //K 
    12'h4c: BcdToAscii = 8'h76; //L 
    12'h4d: BcdToAscii = 8'h77; //M 
    12'h4e: BcdToAscii = 8'h78; //N 
    12'h4f: BcdToAscii = 8'h79; //O 
    12'h50: BcdToAscii = 8'h80; //P 
    12'h51: BcdToAscii = 8'h81; //Q 
    12'h52: BcdToAscii = 8'h82; //R 
    12'h53: BcdToAscii = 8'h83; //S 
    12'h54: BcdToAscii = 8'h84; //T 
    12'h55: BcdToAscii = 8'h85; //U 
    12'h56: BcdToAscii = 8'h86; //V 
    12'h57: BcdToAscii = 8'h87; //W 
    12'h58: BcdToAscii = 8'h88; //X 
    12'h59: BcdToAscii = 8'h89; //Y 
    12'h5a: BcdToAscii = 8'h90; //Z 
    12'h5b: BcdToAscii = 8'h91; //[ 
    12'h5c: BcdToAscii = 8'h92; //\ 
    12'h5d: BcdToAscii = 8'h93; //] 
    12'h5e: BcdToAscii = 8'h94; //^ 
    12'h5f: BcdToAscii = 8'h95; //_ 
    12'h60: BcdToAscii = 8'h96; //` 
    12'h61: BcdToAscii = 8'h97; //a 
    12'h62: BcdToAscii = 8'h98; //b 
    12'h63: BcdToAscii = 8'h99; //c 
    12'h64: BcdToAscii = 8'h100; //d 
    12'h65: BcdToAscii = 8'h101; //e 
    12'h66: BcdToAscii = 8'h102; //f 
    12'h67: BcdToAscii = 8'h103; //g 
    12'h68: BcdToAscii = 8'h104; //h 
    12'h69: BcdToAscii = 8'h105; //i 
    12'h6a: BcdToAscii = 8'h106; //j 
    12'h6b: BcdToAscii = 8'h107; //k 
    12'h6c: BcdToAscii = 8'h108; //l 
    12'h6d: BcdToAscii = 8'h109; //m 
    12'h6e: BcdToAscii = 8'h110; //n 
    12'h6f: BcdToAscii = 8'h111; //o 
    12'h70: BcdToAscii = 8'h112; //p 
    12'h71: BcdToAscii = 8'h113; //q 
    12'h72: BcdToAscii = 8'h114; //r 
    12'h73: BcdToAscii = 8'h115; //s 
    12'h74: BcdToAscii = 8'h116; //t 
    12'h75: BcdToAscii = 8'h117; //u 
    12'h76: BcdToAscii = 8'h118; //v 
    12'h77: BcdToAscii = 8'h119; //w 
    12'h78: BcdToAscii = 8'h120; //x 
    12'h79: BcdToAscii = 8'h121; //y 
    12'h7a: BcdToAscii = 8'h122; //z 
    12'h7b: BcdToAscii = 8'h123; //{ 
    12'h7c: BcdToAscii = 8'h124; //| 
    12'h7d: BcdToAscii = 8'h125; //} 
    12'h7e: BcdToAscii = 8'h126; //~ 
    12'h7f: BcdToAscii = 8'h127; // 
    12'h80: BcdToAscii = 8'h128; // 
    12'h81: BcdToAscii = 8'h129; // 
    12'h82: BcdToAscii = 8'h130; // 
    12'h83: BcdToAscii = 8'h131; // 
    12'h84: BcdToAscii = 8'h132; // 
    12'h85: BcdToAscii = 8'h133; // 
    12'h86: BcdToAscii = 8'h134; // 
    12'h87: BcdToAscii = 8'h135; // 
    12'h88: BcdToAscii = 8'h136; // 
    12'h89: BcdToAscii = 8'h137; // 
    12'h8a: BcdToAscii = 8'h138; // 
    12'h8b: BcdToAscii = 8'h139; // 
    12'h8c: BcdToAscii = 8'h140; // 
    12'h8d: BcdToAscii = 8'h141; // 
    12'h8e: BcdToAscii = 8'h142; // 
    12'h8f: BcdToAscii = 8'h143; // 
    12'h90: BcdToAscii = 8'h144; // 
    12'h91: BcdToAscii = 8'h145; // 
    12'h92: BcdToAscii = 8'h146; // 
    12'h93: BcdToAscii = 8'h147; // 
    12'h94: BcdToAscii = 8'h148; // 
    12'h95: BcdToAscii = 8'h149; // 
    12'h96: BcdToAscii = 8'h150; // 
    12'h97: BcdToAscii = 8'h151; // 
    12'h98: BcdToAscii = 8'h152; // 
    12'h99: BcdToAscii = 8'h153; // 
    12'h9a: BcdToAscii = 8'h154; // 
    12'h9b: BcdToAscii = 8'h155; // 
    12'h9c: BcdToAscii = 8'h156; // 
    12'h9d: BcdToAscii = 8'h157; // 
    12'h9e: BcdToAscii = 8'h158; // 
    12'h9f: BcdToAscii = 8'h159; // 
    12'ha0: BcdToAscii = 8'h160; //  
    12'ha1: BcdToAscii = 8'h161; //¡ 
    12'ha2: BcdToAscii = 8'h162; //¢ 
    12'ha3: BcdToAscii = 8'h163; //£ 
    12'ha4: BcdToAscii = 8'h164; //¤ 
    12'ha5: BcdToAscii = 8'h165; //¥ 
    12'ha6: BcdToAscii = 8'h166; //¦ 
    12'ha7: BcdToAscii = 8'h167; //§ 
    12'ha8: BcdToAscii = 8'h168; //¨ 
    12'ha9: BcdToAscii = 8'h169; //© 
    12'haa: BcdToAscii = 8'h170; //ª 
    12'hab: BcdToAscii = 8'h171; //« 
    12'hac: BcdToAscii = 8'h172; //¬ 
    12'had: BcdToAscii = 8'h173; //­ 
    12'hae: BcdToAscii = 8'h174; //® 
    12'haf: BcdToAscii = 8'h175; //¯ 
    12'hb0: BcdToAscii = 8'h176; //° 
    12'hb1: BcdToAscii = 8'h177; //± 
    12'hb2: BcdToAscii = 8'h178; //² 
    12'hb3: BcdToAscii = 8'h179; //³ 
    12'hb4: BcdToAscii = 8'h180; //´ 
    12'hb5: BcdToAscii = 8'h181; //µ 
    12'hb6: BcdToAscii = 8'h182; //¶ 
    12'hb7: BcdToAscii = 8'h183; //· 
    12'hb8: BcdToAscii = 8'h184; //¸ 
    12'hb9: BcdToAscii = 8'h185; //¹ 
    12'hba: BcdToAscii = 8'h186; //º 
    12'hbb: BcdToAscii = 8'h187; //» 
    12'hbc: BcdToAscii = 8'h188; //¼ 
    12'hbd: BcdToAscii = 8'h189; //½ 
    12'hbe: BcdToAscii = 8'h190; //¾ 
    12'hbf: BcdToAscii = 8'h191; //¿ 
    12'hc0: BcdToAscii = 8'h192; //À 
    12'hc1: BcdToAscii = 8'h193; //Á 
    12'hc2: BcdToAscii = 8'h194; //Â 
    12'hc3: BcdToAscii = 8'h195; //Ã 
    12'hc4: BcdToAscii = 8'h196; //Ä 
    12'hc5: BcdToAscii = 8'h197; //Å 
    12'hc6: BcdToAscii = 8'h198; //Æ 
    12'hc7: BcdToAscii = 8'h199; //Ç 
    12'hc8: BcdToAscii = 8'h200; //È 
    12'hc9: BcdToAscii = 8'h201; //É 
    12'hca: BcdToAscii = 8'h202; //Ê 
    12'hcb: BcdToAscii = 8'h203; //Ë 
    12'hcc: BcdToAscii = 8'h204; //Ì 
    12'hcd: BcdToAscii = 8'h205; //Í 
    12'hce: BcdToAscii = 8'h206; //Î 
    12'hcf: BcdToAscii = 8'h207; //Ï 
    12'hd0: BcdToAscii = 8'h208; //Ð 
    12'hd1: BcdToAscii = 8'h209; //Ñ 
    12'hd2: BcdToAscii = 8'h210; //Ò 
    12'hd3: BcdToAscii = 8'h211; //Ó 
    12'hd4: BcdToAscii = 8'h212; //Ô 
    12'hd5: BcdToAscii = 8'h213; //Õ 
    12'hd6: BcdToAscii = 8'h214; //Ö 
    12'hd7: BcdToAscii = 8'h215; //× 
    12'hd8: BcdToAscii = 8'h216; //Ø 
    12'hd9: BcdToAscii = 8'h217; //Ù 
    12'hda: BcdToAscii = 8'h218; //Ú 
    12'hdb: BcdToAscii = 8'h219; //Û 
    12'hdc: BcdToAscii = 8'h220; //Ü 
    12'hdd: BcdToAscii = 8'h221; //Ý 
    12'hde: BcdToAscii = 8'h222; //Þ 
    12'hdf: BcdToAscii = 8'h223; //ß 
    12'he0: BcdToAscii = 8'h224; //à 
    12'he1: BcdToAscii = 8'h225; //á 
    12'he2: BcdToAscii = 8'h226; //â 
    12'he3: BcdToAscii = 8'h227; //ã 
    12'he4: BcdToAscii = 8'h228; //ä 
    12'he5: BcdToAscii = 8'h229; //å 
    12'he6: BcdToAscii = 8'h230; //æ 
    12'he7: BcdToAscii = 8'h231; //ç 
    12'he8: BcdToAscii = 8'h232; //è 
    12'he9: BcdToAscii = 8'h233; //é 
    12'hea: BcdToAscii = 8'h234; //ê 
    12'heb: BcdToAscii = 8'h235; //ë 
    12'hec: BcdToAscii = 8'h236; //ì 
    12'hed: BcdToAscii = 8'h237; //í 
    12'hee: BcdToAscii = 8'h238; //î 
    12'hef: BcdToAscii = 8'h239; //ï 
    12'hf0: BcdToAscii = 8'h240; //ð 
    12'hf1: BcdToAscii = 8'h241; //ñ 
    12'hf2: BcdToAscii = 8'h242; //ò 
    12'hf3: BcdToAscii = 8'h243; //ó 
    12'hf4: BcdToAscii = 8'h244; //ô 
    12'hf5: BcdToAscii = 8'h245; //õ 
    12'hf6: BcdToAscii = 8'h246; //ö 
    12'hf7: BcdToAscii = 8'h247; //÷ 
    12'hf8: BcdToAscii = 8'h248; //ø 
    12'hf9: BcdToAscii = 8'h249; //ù 
    12'hfa: BcdToAscii = 8'h250; //ú 
    12'hfb: BcdToAscii = 8'h251; //û 
    12'hfc: BcdToAscii = 8'h252; //ü 
    12'hfd: BcdToAscii = 8'h253; //ý 
    12'hfe: BcdToAscii = 8'h254; //þ 
    12'hff: BcdToAscii = 8'h255; //ÿ 
    default: BcdToAscii = {8'bx};n  endcase
endfunction
