`ifndef KEYS_VALUES
   `define KEYS_VALUES

typedef enum  bit [5:0] {
    KEYBOARD_IRAM_KEY =  6'd15,
    KEYBOARD_DRAM_KEY =  6'd10,
    //KEYBOARD_CIN_KEY =  6'd5,
    KEYBOARD_CIO_KEY =  6'd0,

    KEYBOARD_IP_KEY =   6'd35,
    KEYBOARD_LOOP_KEY =  6'd30,
    KEYBOARD_AP_KEY =   6'd25,
    KEYBOARD_DATA_KEY =  6'd20,

    KEYBOARD_0_KEY =    6'd16,
    KEYBOARD_1_KEY =    6'd17,
    KEYBOARD_2_KEY =    6'd18,
    KEYBOARD_3_KEY =    6'd19,
    KEYBOARD_4_KEY =    6'd11,
    KEYBOARD_5_KEY =    6'd12,
    KEYBOARD_6_KEY =    6'd13,
    KEYBOARD_7_KEY =    6'd14,
    KEYBOARD_8_KEY =    6'd6,
    KEYBOARD_9_KEY =    6'd7,
    KEYBOARD_A_KEY =    6'd8,
    KEYBOARD_B_KEY =    6'd9,
    KEYBOARD_C_KEY =    6'd1,
    KEYBOARD_D_KEY =    6'd2,
    KEYBOARD_E_KEY =    6'd3,
    KEYBOARD_F_KEY =    6'd4,

    KEYBOARD_INC_KEY =  6'd36,
    KEYBOARD_DEC_KEY =  6'd31,

    KEYBOARD_HALT_KEY =  6'd26,
    KEYBOARD_STEP_KEY =  6'd33,
    KEYBOARD_RUN_KEY =  6'd28,

    KEYBOARD_ARROW_UP_KEY  =  6'd27,
    KEYBOARD_ARROW_DOWN_KEY = 6'd22,
    KEYBOARD_ARROW_LEFT_KEY = 6'd21,
    KEYBOARD_ARROW_RIGHT_KEY = 6'd23,

    KEYBOARD_HARD_RST =   6'd37,
    KEYBOARD_SOFT_RST_KEY  = 6'd38,

    KEYBOARD_NONAME_KEY =  6'd32,

    KEYBOARD_NONEXIST_2 =  6'd24,
    KEYBOARD_NONEXIST_3 =  6'd29,
    KEYBOARD_NONEXIST_4 =  6'd34
} key_t;

`endif
