`ifndef KEYS_VALUES
   `define KEYS_VALUES

typedef enum   {
    KEYBOARD_IRAM_KEY =  0,
    KEYBOARD_DRAM_KEY =  1,
    KEYBOARD_CIN_KEY =  2,
    KEYBOARD_COUT_KEY =  3,

    KEYBOARD_IP_KEY =   4,
    KEYBOARD_LOOP_KEY =  5,
    KEYBOARD_AP_KEY =   6,
    KEYBOARD_DATA_KEY =  7,

    KEYBOARD_0_KEY =    8,
    KEYBOARD_1_KEY =    16,
    KEYBOARD_2_KEY =    24,
    KEYBOARD_3_KEY =    32,
    KEYBOARD_4_KEY =    9,
    KEYBOARD_5_KEY =    17,
    KEYBOARD_6_KEY =    25,
    KEYBOARD_7_KEY =    33,
    KEYBOARD_8_KEY =    10,
    KEYBOARD_9_KEY =    18,
    KEYBOARD_A_KEY =    26,
    KEYBOARD_B_KEY =    34,
    KEYBOARD_C_KEY =    11,
    KEYBOARD_D_KEY =    19,
    KEYBOARD_E_KEY =    27,
    KEYBOARD_F_KEY =    35,

    KEYBOARD_INC_KEY =  12,
    KEYBOARD_DEC_KEY =  13,

    KEYBOARD_HALT_KEY =  14,
    KEYBOARD_STEP_KEY =  29,
    KEYBOARD_RUN_KEY =  30,

    KEYBOARD_ARROW_UP_KEY  =  22,
    KEYBOARD_ARROW_DOWN_KEY = 23,
    KEYBOARD_ARROW_LEFT_KEY = 15,
    KEYBOARD_ARROW_RIGHT_KEY = 31,

    KEYBOARD_HARD_RST =   20,
    KEYBOARD_SOFT_RST_KEY  = 28,

    KEYBOARD_NONAME_KEY =  21,

    KEYBOARD_NONEXIST_1 =  36,
    KEYBOARD_NONEXIST_2 =  37,
    KEYBOARD_NONEXIST_3 =  38,
    KEYBOARD_NONEXIST_4 =  39
} key_t;

`endif