module ADDSUB(CLOCK, RST, SEQUENCE, ADD, SUB)

parameter SEQUENCE_WIDTH 15

input wire CLOCK;
input wire RST;
input wire[SEQUENCE_WIDTH:0] SEQUENCE;
input wire ADD;
input wire SUB;

always

endmodule
