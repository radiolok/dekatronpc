module dekatronPulseAllow(
    input wire Rst_n,
    input wire Clk,
    input wire En,
    input wire CarryLow,
    input wire CarryHigh,
    //Input pulses:
    input wire [1:0] PulsesIn,
    //Output pulses:
    output wire [1:0] PulsesOut    
);



endmodule