module firmware #(
///home/radiolok/dekatronpc/vhdl/programs/pi/pi.bfk
parameter portSize = 11,
parameter dataSize = 4)(
/* verilator lint_off UNUSEDSIGNAL */
input wire [portSize-1:0] Address,
/* verilator lint_on UNUSEDSIGNAL */
output reg [dataSize-1:0] Data
);
always_comb
/* verilator lint_off WIDTHEXPAND */
  case(Address)
    11'h0: Data = 4'h2; //+ 
    11'h1: Data = 4'h2; //+ 
    11'h2: Data = 4'h2; //+ 
    11'h3: Data = 4'h2; //+ 
    11'h4: Data = 4'h6; //[ 
    11'h5: Data = 4'h5; //< 
    11'h6: Data = 4'h2; //+ 
    11'h7: Data = 4'h4; //> 
    11'h8: Data = 4'h4; //> 
    11'h9: Data = 4'h4; //> 
    11'h10: Data = 4'h4; //> 
    11'h11: Data = 4'h4; //> 
    11'h12: Data = 4'h4; //> 
    11'h13: Data = 4'h4; //> 
    11'h14: Data = 4'h4; //> 
    11'h15: Data = 4'h2; //+ 
    11'h16: Data = 4'h2; //+ 
    11'h17: Data = 4'h2; //+ 
    11'h18: Data = 4'h2; //+ 
    11'h19: Data = 4'h2; //+ 
    11'h20: Data = 4'h2; //+ 
    11'h21: Data = 4'h2; //+ 
    11'h22: Data = 4'h2; //+ 
    11'h23: Data = 4'h2; //+ 
    11'h24: Data = 4'h2; //+ 
    11'h25: Data = 4'h5; //< 
    11'h26: Data = 4'h5; //< 
    11'h27: Data = 4'h5; //< 
    11'h28: Data = 4'h5; //< 
    11'h29: Data = 4'h5; //< 
    11'h30: Data = 4'h5; //< 
    11'h31: Data = 4'h5; //< 
    11'h32: Data = 4'h3; //- 
    11'h33: Data = 4'h7; //] 
    11'h34: Data = 4'h4; //> 
    11'h35: Data = 4'h2; //+ 
    11'h36: Data = 4'h2; //+ 
    11'h37: Data = 4'h2; //+ 
    11'h38: Data = 4'h2; //+ 
    11'h39: Data = 4'h2; //+ 
    11'h40: Data = 4'h6; //[ 
    11'h41: Data = 4'h5; //< 
    11'h42: Data = 4'h2; //+ 
    11'h43: Data = 4'h2; //+ 
    11'h44: Data = 4'h2; //+ 
    11'h45: Data = 4'h2; //+ 
    11'h46: Data = 4'h2; //+ 
    11'h47: Data = 4'h2; //+ 
    11'h48: Data = 4'h2; //+ 
    11'h49: Data = 4'h2; //+ 
    11'h50: Data = 4'h2; //+ 
    11'h51: Data = 4'h4; //> 
    11'h52: Data = 4'h3; //- 
    11'h53: Data = 4'h7; //] 
    11'h54: Data = 4'h2; //+ 
    11'h55: Data = 4'h4; //> 
    11'h56: Data = 4'h4; //> 
    11'h57: Data = 4'h4; //> 
    11'h58: Data = 4'h4; //> 
    11'h59: Data = 4'h4; //> 
    11'h60: Data = 4'h4; //> 
    11'h61: Data = 4'h2; //+ 
    11'h62: Data = 4'h6; //[ 
    11'h63: Data = 4'h5; //< 
    11'h64: Data = 4'h5; //< 
    11'h65: Data = 4'h2; //+ 
    11'h66: Data = 4'h2; //+ 
    11'h67: Data = 4'h2; //+ 
    11'h68: Data = 4'h6; //[ 
    11'h69: Data = 4'h4; //> 
    11'h70: Data = 4'h4; //> 
    11'h71: Data = 4'h6; //[ 
    11'h72: Data = 4'h3; //- 
    11'h73: Data = 4'h5; //< 
    11'h74: Data = 4'h7; //] 
    11'h75: Data = 4'h5; //< 
    11'h76: Data = 4'h6; //[ 
    11'h77: Data = 4'h4; //> 
    11'h78: Data = 4'h7; //] 
    11'h79: Data = 4'h5; //< 
    11'h80: Data = 4'h3; //- 
    11'h81: Data = 4'h7; //] 
    11'h82: Data = 4'h4; //> 
    11'h83: Data = 4'h4; //> 
    11'h84: Data = 4'h6; //[ 
    11'h85: Data = 4'h4; //> 
    11'h86: Data = 4'h2; //+ 
    11'h87: Data = 4'h4; //> 
    11'h88: Data = 4'h7; //] 
    11'h89: Data = 4'h5; //< 
    11'h90: Data = 4'h6; //[ 
    11'h91: Data = 4'h5; //< 
    11'h92: Data = 4'h7; //] 
    11'h93: Data = 4'h4; //> 
    11'h94: Data = 4'h7; //] 
    11'h95: Data = 4'h4; //> 
    11'h96: Data = 4'h6; //[ 
    11'h97: Data = 4'h6; //[ 
    11'h98: Data = 4'h3; //- 
    11'h99: Data = 4'h4; //> 
    11'h100: Data = 4'h4; //> 
    11'h101: Data = 4'h4; //> 
    11'h102: Data = 4'h4; //> 
    11'h103: Data = 4'h2; //+ 
    11'h104: Data = 4'h5; //< 
    11'h105: Data = 4'h5; //< 
    11'h106: Data = 4'h5; //< 
    11'h107: Data = 4'h5; //< 
    11'h108: Data = 4'h7; //] 
    11'h109: Data = 4'h4; //> 
    11'h110: Data = 4'h4; //> 
    11'h111: Data = 4'h4; //> 
    11'h112: Data = 4'h2; //+ 
    11'h113: Data = 4'h2; //+ 
    11'h114: Data = 4'h2; //+ 
    11'h115: Data = 4'h4; //> 
    11'h116: Data = 4'h3; //- 
    11'h117: Data = 4'h7; //] 
    11'h118: Data = 4'h5; //< 
    11'h119: Data = 4'h6; //[ 
    11'h120: Data = 4'h5; //< 
    11'h121: Data = 4'h5; //< 
    11'h122: Data = 4'h5; //< 
    11'h123: Data = 4'h5; //< 
    11'h124: Data = 4'h7; //] 
    11'h125: Data = 4'h5; //< 
    11'h126: Data = 4'h5; //< 
    11'h127: Data = 4'h5; //< 
    11'h128: Data = 4'h5; //< 
    11'h129: Data = 4'h5; //< 
    11'h130: Data = 4'h5; //< 
    11'h131: Data = 4'h5; //< 
    11'h132: Data = 4'h5; //< 
    11'h133: Data = 4'h2; //+ 
    11'h134: Data = 4'h6; //[ 
    11'h135: Data = 4'h3; //- 
    11'h136: Data = 4'h4; //> 
    11'h137: Data = 4'h4; //> 
    11'h138: Data = 4'h4; //> 
    11'h139: Data = 4'h4; //> 
    11'h140: Data = 4'h4; //> 
    11'h141: Data = 4'h4; //> 
    11'h142: Data = 4'h4; //> 
    11'h143: Data = 4'h4; //> 
    11'h144: Data = 4'h4; //> 
    11'h145: Data = 4'h4; //> 
    11'h146: Data = 4'h4; //> 
    11'h147: Data = 4'h4; //> 
    11'h148: Data = 4'h6; //[ 
    11'h149: Data = 4'h5; //< 
    11'h150: Data = 4'h2; //+ 
    11'h151: Data = 4'h6; //[ 
    11'h152: Data = 4'h3; //- 
    11'h153: Data = 4'h4; //> 
    11'h154: Data = 4'h4; //> 
    11'h155: Data = 4'h4; //> 
    11'h156: Data = 4'h4; //> 
    11'h157: Data = 4'h2; //+ 
    11'h158: Data = 4'h5; //< 
    11'h159: Data = 4'h5; //< 
    11'h160: Data = 4'h5; //< 
    11'h161: Data = 4'h5; //< 
    11'h162: Data = 4'h7; //] 
    11'h163: Data = 4'h4; //> 
    11'h164: Data = 4'h4; //> 
    11'h165: Data = 4'h4; //> 
    11'h166: Data = 4'h4; //> 
    11'h167: Data = 4'h4; //> 
    11'h168: Data = 4'h7; //] 
    11'h169: Data = 4'h5; //< 
    11'h170: Data = 4'h5; //< 
    11'h171: Data = 4'h5; //< 
    11'h172: Data = 4'h5; //< 
    11'h173: Data = 4'h6; //[ 
    11'h174: Data = 4'h4; //> 
    11'h175: Data = 4'h4; //> 
    11'h176: Data = 4'h4; //> 
    11'h177: Data = 4'h4; //> 
    11'h178: Data = 4'h4; //> 
    11'h179: Data = 4'h6; //[ 
    11'h180: Data = 4'h5; //< 
    11'h181: Data = 4'h5; //< 
    11'h182: Data = 4'h5; //< 
    11'h183: Data = 4'h5; //< 
    11'h184: Data = 4'h2; //+ 
    11'h185: Data = 4'h4; //> 
    11'h186: Data = 4'h4; //> 
    11'h187: Data = 4'h4; //> 
    11'h188: Data = 4'h4; //> 
    11'h189: Data = 4'h3; //- 
    11'h190: Data = 4'h7; //] 
    11'h191: Data = 4'h5; //< 
    11'h192: Data = 4'h5; //< 
    11'h193: Data = 4'h5; //< 
    11'h194: Data = 4'h5; //< 
    11'h195: Data = 4'h5; //< 
    11'h196: Data = 4'h3; //- 
    11'h197: Data = 4'h6; //[ 
    11'h198: Data = 4'h5; //< 
    11'h199: Data = 4'h5; //< 
    11'h200: Data = 4'h2; //+ 
    11'h201: Data = 4'h2; //+ 
    11'h202: Data = 4'h2; //+ 
    11'h203: Data = 4'h2; //+ 
    11'h204: Data = 4'h2; //+ 
    11'h205: Data = 4'h2; //+ 
    11'h206: Data = 4'h2; //+ 
    11'h207: Data = 4'h2; //+ 
    11'h208: Data = 4'h2; //+ 
    11'h209: Data = 4'h2; //+ 
    11'h210: Data = 4'h4; //> 
    11'h211: Data = 4'h4; //> 
    11'h212: Data = 4'h3; //- 
    11'h213: Data = 4'h7; //] 
    11'h214: Data = 4'h4; //> 
    11'h215: Data = 4'h4; //> 
    11'h216: Data = 4'h4; //> 
    11'h217: Data = 4'h6; //[ 
    11'h218: Data = 4'h5; //< 
    11'h219: Data = 4'h5; //< 
    11'h220: Data = 4'h6; //[ 
    11'h221: Data = 4'h5; //< 
    11'h222: Data = 4'h2; //+ 
    11'h223: Data = 4'h5; //< 
    11'h224: Data = 4'h5; //< 
    11'h225: Data = 4'h2; //+ 
    11'h226: Data = 4'h4; //> 
    11'h227: Data = 4'h4; //> 
    11'h228: Data = 4'h4; //> 
    11'h229: Data = 4'h3; //- 
    11'h230: Data = 4'h7; //] 
    11'h231: Data = 4'h5; //< 
    11'h232: Data = 4'h6; //[ 
    11'h233: Data = 4'h4; //> 
    11'h234: Data = 4'h2; //+ 
    11'h235: Data = 4'h5; //< 
    11'h236: Data = 4'h3; //- 
    11'h237: Data = 4'h7; //] 
    11'h238: Data = 4'h5; //< 
    11'h239: Data = 4'h2; //+ 
    11'h240: Data = 4'h2; //+ 
    11'h241: Data = 4'h5; //< 
    11'h242: Data = 4'h5; //< 
    11'h243: Data = 4'h2; //+ 
    11'h244: Data = 4'h4; //> 
    11'h245: Data = 4'h4; //> 
    11'h246: Data = 4'h4; //> 
    11'h247: Data = 4'h4; //> 
    11'h248: Data = 4'h4; //> 
    11'h249: Data = 4'h4; //> 
    11'h250: Data = 4'h3; //- 
    11'h251: Data = 4'h7; //] 
    11'h252: Data = 4'h5; //< 
    11'h253: Data = 4'h5; //< 
    11'h254: Data = 4'h6; //[ 
    11'h255: Data = 4'h3; //- 
    11'h256: Data = 4'h7; //] 
    11'h257: Data = 4'h5; //< 
    11'h258: Data = 4'h5; //< 
    11'h259: Data = 4'h3; //- 
    11'h260: Data = 4'h5; //< 
    11'h261: Data = 4'h6; //[ 
    11'h262: Data = 4'h3; //- 
    11'h263: Data = 4'h4; //> 
    11'h264: Data = 4'h4; //> 
    11'h265: Data = 4'h2; //+ 
    11'h266: Data = 4'h5; //< 
    11'h267: Data = 4'h3; //- 
    11'h268: Data = 4'h6; //[ 
    11'h269: Data = 4'h4; //> 
    11'h270: Data = 4'h4; //> 
    11'h271: Data = 4'h4; //> 
    11'h272: Data = 4'h7; //] 
    11'h273: Data = 4'h4; //> 
    11'h274: Data = 4'h6; //[ 
    11'h275: Data = 4'h6; //[ 
    11'h276: Data = 4'h5; //< 
    11'h277: Data = 4'h2; //+ 
    11'h278: Data = 4'h4; //> 
    11'h279: Data = 4'h3; //- 
    11'h280: Data = 4'h7; //] 
    11'h281: Data = 4'h4; //> 
    11'h282: Data = 4'h2; //+ 
    11'h283: Data = 4'h4; //> 
    11'h284: Data = 4'h4; //> 
    11'h285: Data = 4'h7; //] 
    11'h286: Data = 4'h5; //< 
    11'h287: Data = 4'h5; //< 
    11'h288: Data = 4'h5; //< 
    11'h289: Data = 4'h5; //< 
    11'h290: Data = 4'h5; //< 
    11'h291: Data = 4'h7; //] 
    11'h292: Data = 4'h4; //> 
    11'h293: Data = 4'h6; //[ 
    11'h294: Data = 4'h3; //- 
    11'h295: Data = 4'h7; //] 
    11'h296: Data = 4'h4; //> 
    11'h297: Data = 4'h2; //+ 
    11'h298: Data = 4'h5; //< 
    11'h299: Data = 4'h5; //< 
    11'h300: Data = 4'h5; //< 
    11'h301: Data = 4'h3; //- 
    11'h302: Data = 4'h6; //[ 
    11'h303: Data = 4'h4; //> 
    11'h304: Data = 4'h4; //> 
    11'h305: Data = 4'h2; //+ 
    11'h306: Data = 4'h5; //< 
    11'h307: Data = 4'h5; //< 
    11'h308: Data = 4'h3; //- 
    11'h309: Data = 4'h7; //] 
    11'h310: Data = 4'h5; //< 
    11'h311: Data = 4'h7; //] 
    11'h312: Data = 4'h5; //< 
    11'h313: Data = 4'h5; //< 
    11'h314: Data = 4'h5; //< 
    11'h315: Data = 4'h5; //< 
    11'h316: Data = 4'h2; //+ 
    11'h317: Data = 4'h4; //> 
    11'h318: Data = 4'h4; //> 
    11'h319: Data = 4'h4; //> 
    11'h320: Data = 4'h4; //> 
    11'h321: Data = 4'h4; //> 
    11'h322: Data = 4'h4; //> 
    11'h323: Data = 4'h4; //> 
    11'h324: Data = 4'h4; //> 
    11'h325: Data = 4'h6; //[ 
    11'h326: Data = 4'h3; //- 
    11'h327: Data = 4'h7; //] 
    11'h328: Data = 4'h4; //> 
    11'h329: Data = 4'h6; //[ 
    11'h330: Data = 4'h5; //< 
    11'h331: Data = 4'h5; //< 
    11'h332: Data = 4'h5; //< 
    11'h333: Data = 4'h2; //+ 
    11'h334: Data = 4'h4; //> 
    11'h335: Data = 4'h4; //> 
    11'h336: Data = 4'h4; //> 
    11'h337: Data = 4'h3; //- 
    11'h338: Data = 4'h7; //] 
    11'h339: Data = 4'h5; //< 
    11'h340: Data = 4'h5; //< 
    11'h341: Data = 4'h2; //+ 
    11'h342: Data = 4'h2; //+ 
    11'h343: Data = 4'h2; //+ 
    11'h344: Data = 4'h2; //+ 
    11'h345: Data = 4'h2; //+ 
    11'h346: Data = 4'h2; //+ 
    11'h347: Data = 4'h2; //+ 
    11'h348: Data = 4'h2; //+ 
    11'h349: Data = 4'h2; //+ 
    11'h350: Data = 4'h2; //+ 
    11'h351: Data = 4'h5; //< 
    11'h352: Data = 4'h6; //[ 
    11'h353: Data = 4'h3; //- 
    11'h354: Data = 4'h4; //> 
    11'h355: Data = 4'h4; //> 
    11'h356: Data = 4'h2; //+ 
    11'h357: Data = 4'h5; //< 
    11'h358: Data = 4'h3; //- 
    11'h359: Data = 4'h6; //[ 
    11'h360: Data = 4'h4; //> 
    11'h361: Data = 4'h4; //> 
    11'h362: Data = 4'h4; //> 
    11'h363: Data = 4'h7; //] 
    11'h364: Data = 4'h4; //> 
    11'h365: Data = 4'h6; //[ 
    11'h366: Data = 4'h6; //[ 
    11'h367: Data = 4'h5; //< 
    11'h368: Data = 4'h2; //+ 
    11'h369: Data = 4'h4; //> 
    11'h370: Data = 4'h3; //- 
    11'h371: Data = 4'h7; //] 
    11'h372: Data = 4'h4; //> 
    11'h373: Data = 4'h2; //+ 
    11'h374: Data = 4'h4; //> 
    11'h375: Data = 4'h4; //> 
    11'h376: Data = 4'h7; //] 
    11'h377: Data = 4'h5; //< 
    11'h378: Data = 4'h5; //< 
    11'h379: Data = 4'h5; //< 
    11'h380: Data = 4'h5; //< 
    11'h381: Data = 4'h5; //< 
    11'h382: Data = 4'h7; //] 
    11'h383: Data = 4'h4; //> 
    11'h384: Data = 4'h6; //[ 
    11'h385: Data = 4'h3; //- 
    11'h386: Data = 4'h7; //] 
    11'h387: Data = 4'h4; //> 
    11'h388: Data = 4'h2; //+ 
    11'h389: Data = 4'h4; //> 
    11'h390: Data = 4'h6; //[ 
    11'h391: Data = 4'h5; //< 
    11'h392: Data = 4'h5; //< 
    11'h393: Data = 4'h2; //+ 
    11'h394: Data = 4'h5; //< 
    11'h395: Data = 4'h2; //+ 
    11'h396: Data = 4'h4; //> 
    11'h397: Data = 4'h4; //> 
    11'h398: Data = 4'h4; //> 
    11'h399: Data = 4'h3; //- 
    11'h400: Data = 4'h7; //] 
    11'h401: Data = 4'h5; //< 
    11'h402: Data = 4'h5; //< 
    11'h403: Data = 4'h5; //< 
    11'h404: Data = 4'h5; //< 
    11'h405: Data = 4'h2; //+ 
    11'h406: Data = 4'h5; //< 
    11'h407: Data = 4'h2; //+ 
    11'h408: Data = 4'h4; //> 
    11'h409: Data = 4'h4; //> 
    11'h410: Data = 4'h6; //[ 
    11'h411: Data = 4'h3; //- 
    11'h412: Data = 4'h6; //[ 
    11'h413: Data = 4'h3; //- 
    11'h414: Data = 4'h6; //[ 
    11'h415: Data = 4'h3; //- 
    11'h416: Data = 4'h6; //[ 
    11'h417: Data = 4'h3; //- 
    11'h418: Data = 4'h6; //[ 
    11'h419: Data = 4'h3; //- 
    11'h420: Data = 4'h6; //[ 
    11'h421: Data = 4'h3; //- 
    11'h422: Data = 4'h6; //[ 
    11'h423: Data = 4'h3; //- 
    11'h424: Data = 4'h6; //[ 
    11'h425: Data = 4'h3; //- 
    11'h426: Data = 4'h6; //[ 
    11'h427: Data = 4'h3; //- 
    11'h428: Data = 4'h5; //< 
    11'h429: Data = 4'h3; //- 
    11'h430: Data = 4'h4; //> 
    11'h431: Data = 4'h6; //[ 
    11'h432: Data = 4'h3; //- 
    11'h433: Data = 4'h5; //< 
    11'h434: Data = 4'h2; //+ 
    11'h435: Data = 4'h5; //< 
    11'h436: Data = 4'h3; //- 
    11'h437: Data = 4'h4; //> 
    11'h438: Data = 4'h4; //> 
    11'h439: Data = 4'h7; //] 
    11'h440: Data = 4'h7; //] 
    11'h441: Data = 4'h7; //] 
    11'h442: Data = 4'h7; //] 
    11'h443: Data = 4'h7; //] 
    11'h444: Data = 4'h7; //] 
    11'h445: Data = 4'h7; //] 
    11'h446: Data = 4'h7; //] 
    11'h447: Data = 4'h7; //] 
    11'h448: Data = 4'h7; //] 
    11'h449: Data = 4'h5; //< 
    11'h450: Data = 4'h6; //[ 
    11'h451: Data = 4'h2; //+ 
    11'h452: Data = 4'h2; //+ 
    11'h453: Data = 4'h2; //+ 
    11'h454: Data = 4'h2; //+ 
    11'h455: Data = 4'h2; //+ 
    11'h456: Data = 4'h6; //[ 
    11'h457: Data = 4'h5; //< 
    11'h458: Data = 4'h5; //< 
    11'h459: Data = 4'h5; //< 
    11'h460: Data = 4'h2; //+ 
    11'h461: Data = 4'h2; //+ 
    11'h462: Data = 4'h2; //+ 
    11'h463: Data = 4'h2; //+ 
    11'h464: Data = 4'h2; //+ 
    11'h465: Data = 4'h2; //+ 
    11'h466: Data = 4'h2; //+ 
    11'h467: Data = 4'h2; //+ 
    11'h468: Data = 4'h5; //< 
    11'h469: Data = 4'h2; //+ 
    11'h470: Data = 4'h2; //+ 
    11'h471: Data = 4'h2; //+ 
    11'h472: Data = 4'h2; //+ 
    11'h473: Data = 4'h2; //+ 
    11'h474: Data = 4'h2; //+ 
    11'h475: Data = 4'h2; //+ 
    11'h476: Data = 4'h2; //+ 
    11'h477: Data = 4'h4; //> 
    11'h478: Data = 4'h4; //> 
    11'h479: Data = 4'h4; //> 
    11'h480: Data = 4'h4; //> 
    11'h481: Data = 4'h3; //- 
    11'h482: Data = 4'h7; //] 
    11'h483: Data = 4'h5; //< 
    11'h484: Data = 4'h5; //< 
    11'h485: Data = 4'h5; //< 
    11'h486: Data = 4'h5; //< 
    11'h487: Data = 4'h2; //+ 
    11'h488: Data = 4'h5; //< 
    11'h489: Data = 4'h3; //- 
    11'h490: Data = 4'h4; //> 
    11'h491: Data = 4'h4; //> 
    11'h492: Data = 4'h4; //> 
    11'h493: Data = 4'h4; //> 
    11'h494: Data = 4'h6; //[ 
    11'h495: Data = 4'h4; //> 
    11'h496: Data = 4'h2; //+ 
    11'h497: Data = 4'h5; //< 
    11'h498: Data = 4'h5; //< 
    11'h499: Data = 4'h5; //< 
    11'h500: Data = 4'h2; //+ 
    11'h501: Data = 4'h2; //+ 
    11'h502: Data = 4'h2; //+ 
    11'h503: Data = 4'h2; //+ 
    11'h504: Data = 4'h2; //+ 
    11'h505: Data = 4'h2; //+ 
    11'h506: Data = 4'h2; //+ 
    11'h507: Data = 4'h2; //+ 
    11'h508: Data = 4'h2; //+ 
    11'h509: Data = 4'h5; //< 
    11'h510: Data = 4'h3; //- 
    11'h511: Data = 4'h4; //> 
    11'h512: Data = 4'h4; //> 
    11'h513: Data = 4'h4; //> 
    11'h514: Data = 4'h3; //- 
    11'h515: Data = 4'h7; //] 
    11'h516: Data = 4'h5; //< 
    11'h517: Data = 4'h5; //< 
    11'h518: Data = 4'h5; //< 
    11'h519: Data = 4'h5; //< 
    11'h520: Data = 4'h5; //< 
    11'h521: Data = 4'h6; //[ 
    11'h522: Data = 4'h4; //> 
    11'h523: Data = 4'h4; //> 
    11'h524: Data = 4'h2; //+ 
    11'h525: Data = 4'h5; //< 
    11'h526: Data = 4'h5; //< 
    11'h527: Data = 4'h3; //- 
    11'h528: Data = 4'h7; //] 
    11'h529: Data = 4'h2; //+ 
    11'h530: Data = 4'h5; //< 
    11'h531: Data = 4'h6; //[ 
    11'h532: Data = 4'h3; //- 
    11'h533: Data = 4'h4; //> 
    11'h534: Data = 4'h3; //- 
    11'h535: Data = 4'h5; //< 
    11'h536: Data = 4'h7; //] 
    11'h537: Data = 4'h4; //> 
    11'h538: Data = 4'h6; //[ 
    11'h539: Data = 4'h4; //> 
    11'h540: Data = 4'h4; //> 
    11'h541: Data = 4'h8; //. 
    11'h542: Data = 4'h5; //< 
    11'h543: Data = 4'h5; //< 
    11'h544: Data = 4'h5; //< 
    11'h545: Data = 4'h5; //< 
    11'h546: Data = 4'h6; //[ 
    11'h547: Data = 4'h2; //+ 
    11'h548: Data = 4'h8; //. 
    11'h549: Data = 4'h6; //[ 
    11'h550: Data = 4'h3; //- 
    11'h551: Data = 4'h7; //] 
    11'h552: Data = 4'h7; //] 
    11'h553: Data = 4'h4; //> 
    11'h554: Data = 4'h4; //> 
    11'h555: Data = 4'h3; //- 
    11'h556: Data = 4'h7; //] 
    11'h557: Data = 4'h4; //> 
    11'h558: Data = 4'h6; //[ 
    11'h559: Data = 4'h4; //> 
    11'h560: Data = 4'h4; //> 
    11'h561: Data = 4'h8; //. 
    11'h562: Data = 4'h5; //< 
    11'h563: Data = 4'h5; //< 
    11'h564: Data = 4'h3; //- 
    11'h565: Data = 4'h7; //] 
    11'h566: Data = 4'h4; //> 
    11'h567: Data = 4'h6; //[ 
    11'h568: Data = 4'h3; //- 
    11'h569: Data = 4'h7; //] 
    11'h570: Data = 4'h4; //> 
    11'h571: Data = 4'h6; //[ 
    11'h572: Data = 4'h3; //- 
    11'h573: Data = 4'h7; //] 
    11'h574: Data = 4'h4; //> 
    11'h575: Data = 4'h4; //> 
    11'h576: Data = 4'h4; //> 
    11'h577: Data = 4'h6; //[ 
    11'h578: Data = 4'h4; //> 
    11'h579: Data = 4'h4; //> 
    11'h580: Data = 4'h6; //[ 
    11'h581: Data = 4'h5; //< 
    11'h582: Data = 4'h5; //< 
    11'h583: Data = 4'h5; //< 
    11'h584: Data = 4'h5; //< 
    11'h585: Data = 4'h5; //< 
    11'h586: Data = 4'h5; //< 
    11'h587: Data = 4'h5; //< 
    11'h588: Data = 4'h5; //< 
    11'h589: Data = 4'h2; //+ 
    11'h590: Data = 4'h4; //> 
    11'h591: Data = 4'h4; //> 
    11'h592: Data = 4'h4; //> 
    11'h593: Data = 4'h4; //> 
    11'h594: Data = 4'h4; //> 
    11'h595: Data = 4'h4; //> 
    11'h596: Data = 4'h4; //> 
    11'h597: Data = 4'h4; //> 
    11'h598: Data = 4'h3; //- 
    11'h599: Data = 4'h7; //] 
    11'h600: Data = 4'h5; //< 
    11'h601: Data = 4'h5; //< 
    11'h602: Data = 4'h3; //- 
    11'h603: Data = 4'h7; //] 
    11'h604: Data = 4'h7; //] 
    11'h605: Data = 4'h4; //> 
    11'h606: Data = 4'h4; //> 
    11'h607: Data = 4'h6; //[ 
    11'h608: Data = 4'h3; //- 
    11'h609: Data = 4'h7; //] 
    11'h610: Data = 4'h5; //< 
    11'h611: Data = 4'h5; //< 
    11'h612: Data = 4'h5; //< 
    11'h613: Data = 4'h6; //[ 
    11'h614: Data = 4'h3; //- 
    11'h615: Data = 4'h7; //] 
    11'h616: Data = 4'h5; //< 
    11'h617: Data = 4'h5; //< 
    11'h618: Data = 4'h5; //< 
    11'h619: Data = 4'h5; //< 
    11'h620: Data = 4'h5; //< 
    11'h621: Data = 4'h5; //< 
    11'h622: Data = 4'h5; //< 
    11'h623: Data = 4'h5; //< 
    11'h624: Data = 4'h7; //] 
    11'h625: Data = 4'h2; //+ 
    11'h626: Data = 4'h2; //+ 
    11'h627: Data = 4'h2; //+ 
    11'h628: Data = 4'h2; //+ 
    11'h629: Data = 4'h2; //+ 
    11'h630: Data = 4'h2; //+ 
    11'h631: Data = 4'h2; //+ 
    11'h632: Data = 4'h2; //+ 
    11'h633: Data = 4'h2; //+ 
    11'h634: Data = 4'h2; //+ 
    11'h635: Data = 4'h8; //. 
    11'h636: Data = 4'h1; //H 
    default: Data = {dataSize{1'bx}};
  endcase

/* verilator lint_on WIDTHEXPAND */
endmodule
