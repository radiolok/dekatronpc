module IpBlock();


endmodule