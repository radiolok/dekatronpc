module helloworld(Address, Data);

parameter portSize = 12;
parameter dataSize = 4;

/* verilator lint_off UNUSEDSIGNAL */
input logic [portSize-1:0] Address;
/* verilator lint_on UNUSEDSIGNAL */
output logic [dataSize-1:0] Data;

always_comb
/* verilator lint_off WIDTHEXPAND */
  case(Address)
    12'b0000: Data = {4'b0010}; //+
    12'b0001: Data = {4'b0010}; //+
    12'b0010: Data = {4'b0010}; //+
    12'b0011: Data = {4'b0010}; //+
    12'b0100: Data = {4'b0010}; //+
    12'b0101: Data = {4'b0010}; //+
    12'b0110: Data = {4'b0010}; //+
    12'b0111: Data = {4'b0010}; //+
    12'b1000: Data = {4'b0010}; //+
    12'b1001: Data = {4'b0010}; //+
    12'b00010000: Data = {4'b0110}; //[
    12'b00010001: Data = {4'b0100}; //>
    12'b00010010: Data = {4'b0010}; //+
    12'b00010011: Data = {4'b0010}; //+
    12'b00010100: Data = {4'b0010}; //+
    12'b00010101: Data = {4'b0010}; //+
    12'b00010110: Data = {4'b0010}; //+
    12'b00010111: Data = {4'b0010}; //+
    12'b00011000: Data = {4'b0010}; //+
    12'b00011001: Data = {4'b0100}; //>
    12'b00100000: Data = {4'b0010}; //+
    12'b00100001: Data = {4'b0010}; //+
    12'b00100010: Data = {4'b0010}; //+
    12'b00100011: Data = {4'b0010}; //+
    12'b00100100: Data = {4'b0010}; //+
    12'b00100101: Data = {4'b0010}; //+
    12'b00100110: Data = {4'b0010}; //+
    12'b00100111: Data = {4'b0010}; //+
    12'b00101000: Data = {4'b0010}; //+
    12'b00101001: Data = {4'b0010}; //+
    12'b00110000: Data = {4'b0100}; //>
    12'b00110001: Data = {4'b0010}; //+
    12'b00110010: Data = {4'b0010}; //+
    12'b00110011: Data = {4'b0010}; //+
    12'b00110100: Data = {4'b0100}; //>
    12'b00110101: Data = {4'b0010}; //+
    12'b00110110: Data = {4'b0101}; //<
    12'b00110111: Data = {4'b0101}; //<
    12'b00111000: Data = {4'b0101}; //<
    12'b00111001: Data = {4'b0101}; //<
    12'b01000000: Data = {4'b0011}; //-
    12'b01000001: Data = {4'b0111}; //]
    12'b01000010: Data = {4'b0100}; //>
    12'b01000011: Data = {4'b0010}; //+
    12'b01000100: Data = {4'b0010}; //+
    12'b01000101: Data = {4'b1000}; //.
    12'b01000110: Data = {4'b0100}; //>
    12'b01000111: Data = {4'b0010}; //+
    12'b01001000: Data = {4'b1000}; //.
    12'b01001001: Data = {4'b0010}; //+
    12'b01010000: Data = {4'b0010}; //+
    12'b01010001: Data = {4'b0010}; //+
    12'b01010010: Data = {4'b0010}; //+
    12'b01010011: Data = {4'b0010}; //+
    12'b01010100: Data = {4'b0010}; //+
    12'b01010101: Data = {4'b0010}; //+
    12'b01010110: Data = {4'b1000}; //.
    12'b01010111: Data = {4'b1000}; //.
    12'b01011000: Data = {4'b0010}; //+
    12'b01011001: Data = {4'b0010}; //+
    12'b01100000: Data = {4'b0010}; //+
    12'b01100001: Data = {4'b1000}; //.
    12'b01100010: Data = {4'b0100}; //>
    12'b01100011: Data = {4'b0010}; //+
    12'b01100100: Data = {4'b0010}; //+
    12'b01100101: Data = {4'b1000}; //.
    12'b01100110: Data = {4'b0101}; //<
    12'b01100111: Data = {4'b0101}; //<
    12'b01101000: Data = {4'b0010}; //+
    12'b01101001: Data = {4'b0010}; //+
    12'b01110000: Data = {4'b0010}; //+
    12'b01110001: Data = {4'b0010}; //+
    12'b01110010: Data = {4'b0010}; //+
    12'b01110011: Data = {4'b0010}; //+
    12'b01110100: Data = {4'b0010}; //+
    12'b01110101: Data = {4'b0010}; //+
    12'b01110110: Data = {4'b0010}; //+
    12'b01110111: Data = {4'b0010}; //+
    12'b01111000: Data = {4'b0010}; //+
    12'b01111001: Data = {4'b0010}; //+
    12'b10000000: Data = {4'b0010}; //+
    12'b10000001: Data = {4'b0010}; //+
    12'b10000010: Data = {4'b0010}; //+
    12'b10000011: Data = {4'b1000}; //.
    12'b10000100: Data = {4'b0100}; //>
    12'b10000101: Data = {4'b1000}; //.
    12'b10000110: Data = {4'b0010}; //+
    12'b10000111: Data = {4'b0010}; //+
    12'b10001000: Data = {4'b0010}; //+
    12'b10001001: Data = {4'b1000}; //.
    12'b10010000: Data = {4'b0011}; //-
    12'b10010001: Data = {4'b0011}; //-
    12'b10010010: Data = {4'b0011}; //-
    12'b10010011: Data = {4'b0011}; //-
    12'b10010100: Data = {4'b0011}; //-
    12'b10010101: Data = {4'b0011}; //-
    12'b10010110: Data = {4'b1000}; //.
    12'b10010111: Data = {4'b0011}; //-
    12'b10011000: Data = {4'b0011}; //-
    12'b10011001: Data = {4'b0011}; //-
    12'b000100000000: Data = {4'b0011}; //-
    12'b000100000001: Data = {4'b0011}; //-
    12'b000100000010: Data = {4'b0011}; //-
    12'b000100000011: Data = {4'b0011}; //-
    12'b000100000100: Data = {4'b0011}; //-
    12'b000100000101: Data = {4'b1000}; //.
    12'b000100000110: Data = {4'b0100}; //>
    12'b000100000111: Data = {4'b0010}; //+
    12'b000100001000: Data = {4'b1000}; //.
    12'b000100001001: Data = {4'b0100}; //>
    12'b000100010000: Data = {4'b1000}; //.
    12'b000100010001: Data = {4'b0001}; //H
    default: Data = {dataSize{1'b0}};
  endcase

/* verilator lint_on WIDTHEXPAND */
endmodule
