module firmware #(
///mnt/d/radiolok@oc.urlnn.ru/Projects/20180271-DekatronPC/vhdl/programs/pi/pi.bfk
parameter portSize = 18,
parameter dataSize = 4)(
/* verilator lint_off UNUSEDSIGNAL */
input wire [portSize-1:0] Address,
/* verilator lint_on UNUSEDSIGNAL */
output reg [dataSize-1:0] Data
);
always_comb
/* verilator lint_off WIDTHEXPAND */
  case(Address)
    18'h0: Data = 4'h2; //+ 
    18'h1: Data = 4'h2; //+ 
    18'h2: Data = 4'h2; //+ 
    18'h3: Data = 4'h2; //+ 
    18'h4: Data = 4'h6; //[ 
    18'h5: Data = 4'h5; //< 
    18'h6: Data = 4'h2; //+ 
    18'h7: Data = 4'h4; //> 
    18'h8: Data = 4'h4; //> 
    18'h9: Data = 4'h4; //> 
    18'h10: Data = 4'h4; //> 
    18'h11: Data = 4'h4; //> 
    18'h12: Data = 4'h4; //> 
    18'h13: Data = 4'h4; //> 
    18'h14: Data = 4'h4; //> 
    18'h15: Data = 4'h2; //+ 
    18'h16: Data = 4'h2; //+ 
    18'h17: Data = 4'h2; //+ 
    18'h18: Data = 4'h2; //+ 
    18'h19: Data = 4'h2; //+ 
    18'h20: Data = 4'h2; //+ 
    18'h21: Data = 4'h2; //+ 
    18'h22: Data = 4'h2; //+ 
    18'h23: Data = 4'h2; //+ 
    18'h24: Data = 4'h2; //+ 
    18'h25: Data = 4'h5; //< 
    18'h26: Data = 4'h5; //< 
    18'h27: Data = 4'h5; //< 
    18'h28: Data = 4'h5; //< 
    18'h29: Data = 4'h5; //< 
    18'h30: Data = 4'h5; //< 
    18'h31: Data = 4'h5; //< 
    18'h32: Data = 4'h3; //- 
    18'h33: Data = 4'h7; //] 
    18'h34: Data = 4'h4; //> 
    18'h35: Data = 4'h2; //+ 
    18'h36: Data = 4'h2; //+ 
    18'h37: Data = 4'h2; //+ 
    18'h38: Data = 4'h2; //+ 
    18'h39: Data = 4'h2; //+ 
    18'h40: Data = 4'h6; //[ 
    18'h41: Data = 4'h5; //< 
    18'h42: Data = 4'h2; //+ 
    18'h43: Data = 4'h2; //+ 
    18'h44: Data = 4'h2; //+ 
    18'h45: Data = 4'h2; //+ 
    18'h46: Data = 4'h2; //+ 
    18'h47: Data = 4'h2; //+ 
    18'h48: Data = 4'h2; //+ 
    18'h49: Data = 4'h2; //+ 
    18'h50: Data = 4'h2; //+ 
    18'h51: Data = 4'h4; //> 
    18'h52: Data = 4'h3; //- 
    18'h53: Data = 4'h7; //] 
    18'h54: Data = 4'h2; //+ 
    18'h55: Data = 4'h4; //> 
    18'h56: Data = 4'h4; //> 
    18'h57: Data = 4'h4; //> 
    18'h58: Data = 4'h4; //> 
    18'h59: Data = 4'h4; //> 
    18'h60: Data = 4'h4; //> 
    18'h61: Data = 4'h2; //+ 
    18'h62: Data = 4'h6; //[ 
    18'h63: Data = 4'h5; //< 
    18'h64: Data = 4'h5; //< 
    18'h65: Data = 4'h2; //+ 
    18'h66: Data = 4'h2; //+ 
    18'h67: Data = 4'h2; //+ 
    18'h68: Data = 4'h6; //[ 
    18'h69: Data = 4'h4; //> 
    18'h70: Data = 4'h4; //> 
    18'h71: Data = 4'h6; //[ 
    18'h72: Data = 4'h3; //- 
    18'h73: Data = 4'h5; //< 
    18'h74: Data = 4'h7; //] 
    18'h75: Data = 4'h5; //< 
    18'h76: Data = 4'h6; //[ 
    18'h77: Data = 4'h4; //> 
    18'h78: Data = 4'h7; //] 
    18'h79: Data = 4'h5; //< 
    18'h80: Data = 4'h3; //- 
    18'h81: Data = 4'h7; //] 
    18'h82: Data = 4'h4; //> 
    18'h83: Data = 4'h4; //> 
    18'h84: Data = 4'h6; //[ 
    18'h85: Data = 4'h4; //> 
    18'h86: Data = 4'h2; //+ 
    18'h87: Data = 4'h4; //> 
    18'h88: Data = 4'h7; //] 
    18'h89: Data = 4'h5; //< 
    18'h90: Data = 4'h6; //[ 
    18'h91: Data = 4'h5; //< 
    18'h92: Data = 4'h7; //] 
    18'h93: Data = 4'h4; //> 
    18'h94: Data = 4'h7; //] 
    18'h95: Data = 4'h4; //> 
    18'h96: Data = 4'h6; //[ 
    18'h97: Data = 4'h6; //[ 
    18'h98: Data = 4'h3; //- 
    18'h99: Data = 4'h4; //> 
    18'h100: Data = 4'h4; //> 
    18'h101: Data = 4'h4; //> 
    18'h102: Data = 4'h4; //> 
    18'h103: Data = 4'h2; //+ 
    18'h104: Data = 4'h5; //< 
    18'h105: Data = 4'h5; //< 
    18'h106: Data = 4'h5; //< 
    18'h107: Data = 4'h5; //< 
    18'h108: Data = 4'h7; //] 
    18'h109: Data = 4'h4; //> 
    18'h110: Data = 4'h4; //> 
    18'h111: Data = 4'h4; //> 
    18'h112: Data = 4'h2; //+ 
    18'h113: Data = 4'h2; //+ 
    18'h114: Data = 4'h2; //+ 
    18'h115: Data = 4'h4; //> 
    18'h116: Data = 4'h3; //- 
    18'h117: Data = 4'h7; //] 
    18'h118: Data = 4'h5; //< 
    18'h119: Data = 4'h6; //[ 
    18'h120: Data = 4'h5; //< 
    18'h121: Data = 4'h5; //< 
    18'h122: Data = 4'h5; //< 
    18'h123: Data = 4'h5; //< 
    18'h124: Data = 4'h7; //] 
    18'h125: Data = 4'h5; //< 
    18'h126: Data = 4'h5; //< 
    18'h127: Data = 4'h5; //< 
    18'h128: Data = 4'h5; //< 
    18'h129: Data = 4'h5; //< 
    18'h130: Data = 4'h5; //< 
    18'h131: Data = 4'h5; //< 
    18'h132: Data = 4'h5; //< 
    18'h133: Data = 4'h2; //+ 
    18'h134: Data = 4'h6; //[ 
    18'h135: Data = 4'h3; //- 
    18'h136: Data = 4'h4; //> 
    18'h137: Data = 4'h4; //> 
    18'h138: Data = 4'h4; //> 
    18'h139: Data = 4'h4; //> 
    18'h140: Data = 4'h4; //> 
    18'h141: Data = 4'h4; //> 
    18'h142: Data = 4'h4; //> 
    18'h143: Data = 4'h4; //> 
    18'h144: Data = 4'h4; //> 
    18'h145: Data = 4'h4; //> 
    18'h146: Data = 4'h4; //> 
    18'h147: Data = 4'h4; //> 
    18'h148: Data = 4'h6; //[ 
    18'h149: Data = 4'h5; //< 
    18'h150: Data = 4'h2; //+ 
    18'h151: Data = 4'h6; //[ 
    18'h152: Data = 4'h3; //- 
    18'h153: Data = 4'h4; //> 
    18'h154: Data = 4'h4; //> 
    18'h155: Data = 4'h4; //> 
    18'h156: Data = 4'h4; //> 
    18'h157: Data = 4'h2; //+ 
    18'h158: Data = 4'h5; //< 
    18'h159: Data = 4'h5; //< 
    18'h160: Data = 4'h5; //< 
    18'h161: Data = 4'h5; //< 
    18'h162: Data = 4'h7; //] 
    18'h163: Data = 4'h4; //> 
    18'h164: Data = 4'h4; //> 
    18'h165: Data = 4'h4; //> 
    18'h166: Data = 4'h4; //> 
    18'h167: Data = 4'h4; //> 
    18'h168: Data = 4'h7; //] 
    18'h169: Data = 4'h5; //< 
    18'h170: Data = 4'h5; //< 
    18'h171: Data = 4'h5; //< 
    18'h172: Data = 4'h5; //< 
    18'h173: Data = 4'h6; //[ 
    18'h174: Data = 4'h4; //> 
    18'h175: Data = 4'h4; //> 
    18'h176: Data = 4'h4; //> 
    18'h177: Data = 4'h4; //> 
    18'h178: Data = 4'h4; //> 
    18'h179: Data = 4'h6; //[ 
    18'h180: Data = 4'h5; //< 
    18'h181: Data = 4'h5; //< 
    18'h182: Data = 4'h5; //< 
    18'h183: Data = 4'h5; //< 
    18'h184: Data = 4'h2; //+ 
    18'h185: Data = 4'h4; //> 
    18'h186: Data = 4'h4; //> 
    18'h187: Data = 4'h4; //> 
    18'h188: Data = 4'h4; //> 
    18'h189: Data = 4'h3; //- 
    18'h190: Data = 4'h7; //] 
    18'h191: Data = 4'h5; //< 
    18'h192: Data = 4'h5; //< 
    18'h193: Data = 4'h5; //< 
    18'h194: Data = 4'h5; //< 
    18'h195: Data = 4'h5; //< 
    18'h196: Data = 4'h3; //- 
    18'h197: Data = 4'h6; //[ 
    18'h198: Data = 4'h5; //< 
    18'h199: Data = 4'h5; //< 
    18'h200: Data = 4'h2; //+ 
    18'h201: Data = 4'h2; //+ 
    18'h202: Data = 4'h2; //+ 
    18'h203: Data = 4'h2; //+ 
    18'h204: Data = 4'h2; //+ 
    18'h205: Data = 4'h2; //+ 
    18'h206: Data = 4'h2; //+ 
    18'h207: Data = 4'h2; //+ 
    18'h208: Data = 4'h2; //+ 
    18'h209: Data = 4'h2; //+ 
    18'h210: Data = 4'h4; //> 
    18'h211: Data = 4'h4; //> 
    18'h212: Data = 4'h3; //- 
    18'h213: Data = 4'h7; //] 
    18'h214: Data = 4'h4; //> 
    18'h215: Data = 4'h4; //> 
    18'h216: Data = 4'h4; //> 
    18'h217: Data = 4'h6; //[ 
    18'h218: Data = 4'h5; //< 
    18'h219: Data = 4'h5; //< 
    18'h220: Data = 4'h6; //[ 
    18'h221: Data = 4'h5; //< 
    18'h222: Data = 4'h2; //+ 
    18'h223: Data = 4'h5; //< 
    18'h224: Data = 4'h5; //< 
    18'h225: Data = 4'h2; //+ 
    18'h226: Data = 4'h4; //> 
    18'h227: Data = 4'h4; //> 
    18'h228: Data = 4'h4; //> 
    18'h229: Data = 4'h3; //- 
    18'h230: Data = 4'h7; //] 
    18'h231: Data = 4'h5; //< 
    18'h232: Data = 4'h6; //[ 
    18'h233: Data = 4'h4; //> 
    18'h234: Data = 4'h2; //+ 
    18'h235: Data = 4'h5; //< 
    18'h236: Data = 4'h3; //- 
    18'h237: Data = 4'h7; //] 
    18'h238: Data = 4'h5; //< 
    18'h239: Data = 4'h2; //+ 
    18'h240: Data = 4'h2; //+ 
    18'h241: Data = 4'h5; //< 
    18'h242: Data = 4'h5; //< 
    18'h243: Data = 4'h2; //+ 
    18'h244: Data = 4'h4; //> 
    18'h245: Data = 4'h4; //> 
    18'h246: Data = 4'h4; //> 
    18'h247: Data = 4'h4; //> 
    18'h248: Data = 4'h4; //> 
    18'h249: Data = 4'h4; //> 
    18'h250: Data = 4'h3; //- 
    18'h251: Data = 4'h7; //] 
    18'h252: Data = 4'h5; //< 
    18'h253: Data = 4'h5; //< 
    18'h254: Data = 4'h6; //[ 
    18'h255: Data = 4'h3; //- 
    18'h256: Data = 4'h7; //] 
    18'h257: Data = 4'h5; //< 
    18'h258: Data = 4'h5; //< 
    18'h259: Data = 4'h3; //- 
    18'h260: Data = 4'h5; //< 
    18'h261: Data = 4'h6; //[ 
    18'h262: Data = 4'h3; //- 
    18'h263: Data = 4'h4; //> 
    18'h264: Data = 4'h4; //> 
    18'h265: Data = 4'h2; //+ 
    18'h266: Data = 4'h5; //< 
    18'h267: Data = 4'h3; //- 
    18'h268: Data = 4'h6; //[ 
    18'h269: Data = 4'h4; //> 
    18'h270: Data = 4'h4; //> 
    18'h271: Data = 4'h4; //> 
    18'h272: Data = 4'h7; //] 
    18'h273: Data = 4'h4; //> 
    18'h274: Data = 4'h6; //[ 
    18'h275: Data = 4'h6; //[ 
    18'h276: Data = 4'h5; //< 
    18'h277: Data = 4'h2; //+ 
    18'h278: Data = 4'h4; //> 
    18'h279: Data = 4'h3; //- 
    18'h280: Data = 4'h7; //] 
    18'h281: Data = 4'h4; //> 
    18'h282: Data = 4'h2; //+ 
    18'h283: Data = 4'h4; //> 
    18'h284: Data = 4'h4; //> 
    18'h285: Data = 4'h7; //] 
    18'h286: Data = 4'h5; //< 
    18'h287: Data = 4'h5; //< 
    18'h288: Data = 4'h5; //< 
    18'h289: Data = 4'h5; //< 
    18'h290: Data = 4'h5; //< 
    18'h291: Data = 4'h7; //] 
    18'h292: Data = 4'h4; //> 
    18'h293: Data = 4'h6; //[ 
    18'h294: Data = 4'h3; //- 
    18'h295: Data = 4'h7; //] 
    18'h296: Data = 4'h4; //> 
    18'h297: Data = 4'h2; //+ 
    18'h298: Data = 4'h5; //< 
    18'h299: Data = 4'h5; //< 
    18'h300: Data = 4'h5; //< 
    18'h301: Data = 4'h3; //- 
    18'h302: Data = 4'h6; //[ 
    18'h303: Data = 4'h4; //> 
    18'h304: Data = 4'h4; //> 
    18'h305: Data = 4'h2; //+ 
    18'h306: Data = 4'h5; //< 
    18'h307: Data = 4'h5; //< 
    18'h308: Data = 4'h3; //- 
    18'h309: Data = 4'h7; //] 
    18'h310: Data = 4'h5; //< 
    18'h311: Data = 4'h7; //] 
    18'h312: Data = 4'h5; //< 
    18'h313: Data = 4'h5; //< 
    18'h314: Data = 4'h5; //< 
    18'h315: Data = 4'h5; //< 
    18'h316: Data = 4'h2; //+ 
    18'h317: Data = 4'h4; //> 
    18'h318: Data = 4'h4; //> 
    18'h319: Data = 4'h4; //> 
    18'h320: Data = 4'h4; //> 
    18'h321: Data = 4'h4; //> 
    18'h322: Data = 4'h4; //> 
    18'h323: Data = 4'h4; //> 
    18'h324: Data = 4'h4; //> 
    18'h325: Data = 4'h6; //[ 
    18'h326: Data = 4'h3; //- 
    18'h327: Data = 4'h7; //] 
    18'h328: Data = 4'h4; //> 
    18'h329: Data = 4'h6; //[ 
    18'h330: Data = 4'h5; //< 
    18'h331: Data = 4'h5; //< 
    18'h332: Data = 4'h5; //< 
    18'h333: Data = 4'h2; //+ 
    18'h334: Data = 4'h4; //> 
    18'h335: Data = 4'h4; //> 
    18'h336: Data = 4'h4; //> 
    18'h337: Data = 4'h3; //- 
    18'h338: Data = 4'h7; //] 
    18'h339: Data = 4'h5; //< 
    18'h340: Data = 4'h5; //< 
    18'h341: Data = 4'h2; //+ 
    18'h342: Data = 4'h2; //+ 
    18'h343: Data = 4'h2; //+ 
    18'h344: Data = 4'h2; //+ 
    18'h345: Data = 4'h2; //+ 
    18'h346: Data = 4'h2; //+ 
    18'h347: Data = 4'h2; //+ 
    18'h348: Data = 4'h2; //+ 
    18'h349: Data = 4'h2; //+ 
    18'h350: Data = 4'h2; //+ 
    18'h351: Data = 4'h5; //< 
    18'h352: Data = 4'h6; //[ 
    18'h353: Data = 4'h3; //- 
    18'h354: Data = 4'h4; //> 
    18'h355: Data = 4'h4; //> 
    18'h356: Data = 4'h2; //+ 
    18'h357: Data = 4'h5; //< 
    18'h358: Data = 4'h3; //- 
    18'h359: Data = 4'h6; //[ 
    18'h360: Data = 4'h4; //> 
    18'h361: Data = 4'h4; //> 
    18'h362: Data = 4'h4; //> 
    18'h363: Data = 4'h7; //] 
    18'h364: Data = 4'h4; //> 
    18'h365: Data = 4'h6; //[ 
    18'h366: Data = 4'h6; //[ 
    18'h367: Data = 4'h5; //< 
    18'h368: Data = 4'h2; //+ 
    18'h369: Data = 4'h4; //> 
    18'h370: Data = 4'h3; //- 
    18'h371: Data = 4'h7; //] 
    18'h372: Data = 4'h4; //> 
    18'h373: Data = 4'h2; //+ 
    18'h374: Data = 4'h4; //> 
    18'h375: Data = 4'h4; //> 
    18'h376: Data = 4'h7; //] 
    18'h377: Data = 4'h5; //< 
    18'h378: Data = 4'h5; //< 
    18'h379: Data = 4'h5; //< 
    18'h380: Data = 4'h5; //< 
    18'h381: Data = 4'h5; //< 
    18'h382: Data = 4'h7; //] 
    18'h383: Data = 4'h4; //> 
    18'h384: Data = 4'h6; //[ 
    18'h385: Data = 4'h3; //- 
    18'h386: Data = 4'h7; //] 
    18'h387: Data = 4'h4; //> 
    18'h388: Data = 4'h2; //+ 
    18'h389: Data = 4'h4; //> 
    18'h390: Data = 4'h6; //[ 
    18'h391: Data = 4'h5; //< 
    18'h392: Data = 4'h5; //< 
    18'h393: Data = 4'h2; //+ 
    18'h394: Data = 4'h5; //< 
    18'h395: Data = 4'h2; //+ 
    18'h396: Data = 4'h4; //> 
    18'h397: Data = 4'h4; //> 
    18'h398: Data = 4'h4; //> 
    18'h399: Data = 4'h3; //- 
    18'h400: Data = 4'h7; //] 
    18'h401: Data = 4'h5; //< 
    18'h402: Data = 4'h5; //< 
    18'h403: Data = 4'h5; //< 
    18'h404: Data = 4'h5; //< 
    18'h405: Data = 4'h2; //+ 
    18'h406: Data = 4'h5; //< 
    18'h407: Data = 4'h2; //+ 
    18'h408: Data = 4'h4; //> 
    18'h409: Data = 4'h4; //> 
    18'h410: Data = 4'h6; //[ 
    18'h411: Data = 4'h3; //- 
    18'h412: Data = 4'h6; //[ 
    18'h413: Data = 4'h3; //- 
    18'h414: Data = 4'h6; //[ 
    18'h415: Data = 4'h3; //- 
    18'h416: Data = 4'h6; //[ 
    18'h417: Data = 4'h3; //- 
    18'h418: Data = 4'h6; //[ 
    18'h419: Data = 4'h3; //- 
    18'h420: Data = 4'h6; //[ 
    18'h421: Data = 4'h3; //- 
    18'h422: Data = 4'h6; //[ 
    18'h423: Data = 4'h3; //- 
    18'h424: Data = 4'h6; //[ 
    18'h425: Data = 4'h3; //- 
    18'h426: Data = 4'h6; //[ 
    18'h427: Data = 4'h3; //- 
    18'h428: Data = 4'h5; //< 
    18'h429: Data = 4'h3; //- 
    18'h430: Data = 4'h4; //> 
    18'h431: Data = 4'h6; //[ 
    18'h432: Data = 4'h3; //- 
    18'h433: Data = 4'h5; //< 
    18'h434: Data = 4'h2; //+ 
    18'h435: Data = 4'h5; //< 
    18'h436: Data = 4'h3; //- 
    18'h437: Data = 4'h4; //> 
    18'h438: Data = 4'h4; //> 
    18'h439: Data = 4'h7; //] 
    18'h440: Data = 4'h7; //] 
    18'h441: Data = 4'h7; //] 
    18'h442: Data = 4'h7; //] 
    18'h443: Data = 4'h7; //] 
    18'h444: Data = 4'h7; //] 
    18'h445: Data = 4'h7; //] 
    18'h446: Data = 4'h7; //] 
    18'h447: Data = 4'h7; //] 
    18'h448: Data = 4'h7; //] 
    18'h449: Data = 4'h5; //< 
    18'h450: Data = 4'h6; //[ 
    18'h451: Data = 4'h2; //+ 
    18'h452: Data = 4'h2; //+ 
    18'h453: Data = 4'h2; //+ 
    18'h454: Data = 4'h2; //+ 
    18'h455: Data = 4'h2; //+ 
    18'h456: Data = 4'h6; //[ 
    18'h457: Data = 4'h5; //< 
    18'h458: Data = 4'h5; //< 
    18'h459: Data = 4'h5; //< 
    18'h460: Data = 4'h2; //+ 
    18'h461: Data = 4'h2; //+ 
    18'h462: Data = 4'h2; //+ 
    18'h463: Data = 4'h2; //+ 
    18'h464: Data = 4'h2; //+ 
    18'h465: Data = 4'h2; //+ 
    18'h466: Data = 4'h2; //+ 
    18'h467: Data = 4'h2; //+ 
    18'h468: Data = 4'h5; //< 
    18'h469: Data = 4'h2; //+ 
    18'h470: Data = 4'h2; //+ 
    18'h471: Data = 4'h2; //+ 
    18'h472: Data = 4'h2; //+ 
    18'h473: Data = 4'h2; //+ 
    18'h474: Data = 4'h2; //+ 
    18'h475: Data = 4'h2; //+ 
    18'h476: Data = 4'h2; //+ 
    18'h477: Data = 4'h4; //> 
    18'h478: Data = 4'h4; //> 
    18'h479: Data = 4'h4; //> 
    18'h480: Data = 4'h4; //> 
    18'h481: Data = 4'h3; //- 
    18'h482: Data = 4'h7; //] 
    18'h483: Data = 4'h5; //< 
    18'h484: Data = 4'h5; //< 
    18'h485: Data = 4'h5; //< 
    18'h486: Data = 4'h5; //< 
    18'h487: Data = 4'h2; //+ 
    18'h488: Data = 4'h5; //< 
    18'h489: Data = 4'h3; //- 
    18'h490: Data = 4'h4; //> 
    18'h491: Data = 4'h4; //> 
    18'h492: Data = 4'h4; //> 
    18'h493: Data = 4'h4; //> 
    18'h494: Data = 4'h6; //[ 
    18'h495: Data = 4'h4; //> 
    18'h496: Data = 4'h2; //+ 
    18'h497: Data = 4'h5; //< 
    18'h498: Data = 4'h5; //< 
    18'h499: Data = 4'h5; //< 
    18'h500: Data = 4'h2; //+ 
    18'h501: Data = 4'h2; //+ 
    18'h502: Data = 4'h2; //+ 
    18'h503: Data = 4'h2; //+ 
    18'h504: Data = 4'h2; //+ 
    18'h505: Data = 4'h2; //+ 
    18'h506: Data = 4'h2; //+ 
    18'h507: Data = 4'h2; //+ 
    18'h508: Data = 4'h2; //+ 
    18'h509: Data = 4'h5; //< 
    18'h510: Data = 4'h3; //- 
    18'h511: Data = 4'h4; //> 
    18'h512: Data = 4'h4; //> 
    18'h513: Data = 4'h4; //> 
    18'h514: Data = 4'h3; //- 
    18'h515: Data = 4'h7; //] 
    18'h516: Data = 4'h5; //< 
    18'h517: Data = 4'h5; //< 
    18'h518: Data = 4'h5; //< 
    18'h519: Data = 4'h5; //< 
    18'h520: Data = 4'h5; //< 
    18'h521: Data = 4'h6; //[ 
    18'h522: Data = 4'h4; //> 
    18'h523: Data = 4'h4; //> 
    18'h524: Data = 4'h2; //+ 
    18'h525: Data = 4'h5; //< 
    18'h526: Data = 4'h5; //< 
    18'h527: Data = 4'h3; //- 
    18'h528: Data = 4'h7; //] 
    18'h529: Data = 4'h2; //+ 
    18'h530: Data = 4'h5; //< 
    18'h531: Data = 4'h6; //[ 
    18'h532: Data = 4'h3; //- 
    18'h533: Data = 4'h4; //> 
    18'h534: Data = 4'h3; //- 
    18'h535: Data = 4'h5; //< 
    18'h536: Data = 4'h7; //] 
    18'h537: Data = 4'h4; //> 
    18'h538: Data = 4'h6; //[ 
    18'h539: Data = 4'h4; //> 
    18'h540: Data = 4'h4; //> 
    18'h541: Data = 4'h8; //. 
    18'h542: Data = 4'h5; //< 
    18'h543: Data = 4'h5; //< 
    18'h544: Data = 4'h5; //< 
    18'h545: Data = 4'h5; //< 
    18'h546: Data = 4'h6; //[ 
    18'h547: Data = 4'h2; //+ 
    18'h548: Data = 4'h8; //. 
    18'h549: Data = 4'h6; //[ 
    18'h550: Data = 4'h3; //- 
    18'h551: Data = 4'h7; //] 
    18'h552: Data = 4'h7; //] 
    18'h553: Data = 4'h4; //> 
    18'h554: Data = 4'h4; //> 
    18'h555: Data = 4'h3; //- 
    18'h556: Data = 4'h7; //] 
    18'h557: Data = 4'h4; //> 
    18'h558: Data = 4'h6; //[ 
    18'h559: Data = 4'h4; //> 
    18'h560: Data = 4'h4; //> 
    18'h561: Data = 4'h8; //. 
    18'h562: Data = 4'h5; //< 
    18'h563: Data = 4'h5; //< 
    18'h564: Data = 4'h3; //- 
    18'h565: Data = 4'h7; //] 
    18'h566: Data = 4'h4; //> 
    18'h567: Data = 4'h6; //[ 
    18'h568: Data = 4'h3; //- 
    18'h569: Data = 4'h7; //] 
    18'h570: Data = 4'h4; //> 
    18'h571: Data = 4'h6; //[ 
    18'h572: Data = 4'h3; //- 
    18'h573: Data = 4'h7; //] 
    18'h574: Data = 4'h4; //> 
    18'h575: Data = 4'h4; //> 
    18'h576: Data = 4'h4; //> 
    18'h577: Data = 4'h6; //[ 
    18'h578: Data = 4'h4; //> 
    18'h579: Data = 4'h4; //> 
    18'h580: Data = 4'h6; //[ 
    18'h581: Data = 4'h5; //< 
    18'h582: Data = 4'h5; //< 
    18'h583: Data = 4'h5; //< 
    18'h584: Data = 4'h5; //< 
    18'h585: Data = 4'h5; //< 
    18'h586: Data = 4'h5; //< 
    18'h587: Data = 4'h5; //< 
    18'h588: Data = 4'h5; //< 
    18'h589: Data = 4'h2; //+ 
    18'h590: Data = 4'h4; //> 
    18'h591: Data = 4'h4; //> 
    18'h592: Data = 4'h4; //> 
    18'h593: Data = 4'h4; //> 
    18'h594: Data = 4'h4; //> 
    18'h595: Data = 4'h4; //> 
    18'h596: Data = 4'h4; //> 
    18'h597: Data = 4'h4; //> 
    18'h598: Data = 4'h3; //- 
    18'h599: Data = 4'h7; //] 
    18'h600: Data = 4'h5; //< 
    18'h601: Data = 4'h5; //< 
    18'h602: Data = 4'h3; //- 
    18'h603: Data = 4'h7; //] 
    18'h604: Data = 4'h7; //] 
    18'h605: Data = 4'h4; //> 
    18'h606: Data = 4'h4; //> 
    18'h607: Data = 4'h6; //[ 
    18'h608: Data = 4'h3; //- 
    18'h609: Data = 4'h7; //] 
    18'h610: Data = 4'h5; //< 
    18'h611: Data = 4'h5; //< 
    18'h612: Data = 4'h5; //< 
    18'h613: Data = 4'h6; //[ 
    18'h614: Data = 4'h3; //- 
    18'h615: Data = 4'h7; //] 
    18'h616: Data = 4'h5; //< 
    18'h617: Data = 4'h5; //< 
    18'h618: Data = 4'h5; //< 
    18'h619: Data = 4'h5; //< 
    18'h620: Data = 4'h5; //< 
    18'h621: Data = 4'h5; //< 
    18'h622: Data = 4'h5; //< 
    18'h623: Data = 4'h5; //< 
    18'h624: Data = 4'h7; //] 
    18'h625: Data = 4'h2; //+ 
    18'h626: Data = 4'h2; //+ 
    18'h627: Data = 4'h2; //+ 
    18'h628: Data = 4'h2; //+ 
    18'h629: Data = 4'h2; //+ 
    18'h630: Data = 4'h2; //+ 
    18'h631: Data = 4'h2; //+ 
    18'h632: Data = 4'h2; //+ 
    18'h633: Data = 4'h2; //+ 
    18'h634: Data = 4'h2; //+ 
    18'h635: Data = 4'h8; //. 
    18'h636: Data = 4'h1; //H 
    18'h10000: Data = 4'h2; //+ 
    18'h10001: Data = 4'h2; //+ 
    18'h10002: Data = 4'h2; //+ 
    18'h10003: Data = 4'h2; //+ 
    18'h10004: Data = 4'h2; //+ 
    18'h10005: Data = 4'h2; //+ 
    18'h10006: Data = 4'h2; //+ 
    18'h10007: Data = 4'h2; //+ 
    18'h10008: Data = 4'h2; //+ 
    18'h10009: Data = 4'h2; //+ 
    18'h10010: Data = 4'h2; //+ 
    18'h10011: Data = 4'h2; //+ 
    18'h10012: Data = 4'h2; //+ 
    18'h10013: Data = 4'h6; //[ 
    18'h10014: Data = 4'h3; //- 
    18'h10015: Data = 4'h4; //> 
    18'h10016: Data = 4'h2; //+ 
    18'h10017: Data = 4'h2; //+ 
    18'h10018: Data = 4'h4; //> 
    18'h10019: Data = 4'h4; //> 
    18'h10020: Data = 4'h4; //> 
    18'h10021: Data = 4'h2; //+ 
    18'h10022: Data = 4'h2; //+ 
    18'h10023: Data = 4'h2; //+ 
    18'h10024: Data = 4'h2; //+ 
    18'h10025: Data = 4'h2; //+ 
    18'h10026: Data = 4'h4; //> 
    18'h10027: Data = 4'h2; //+ 
    18'h10028: Data = 4'h2; //+ 
    18'h10029: Data = 4'h4; //> 
    18'h10030: Data = 4'h2; //+ 
    18'h10031: Data = 4'h5; //< 
    18'h10032: Data = 4'h5; //< 
    18'h10033: Data = 4'h5; //< 
    18'h10034: Data = 4'h5; //< 
    18'h10035: Data = 4'h5; //< 
    18'h10036: Data = 4'h5; //< 
    18'h10037: Data = 4'h7; //] 
    18'h10038: Data = 4'h4; //> 
    18'h10039: Data = 4'h4; //> 
    18'h10040: Data = 4'h4; //> 
    18'h10041: Data = 4'h4; //> 
    18'h10042: Data = 4'h4; //> 
    18'h10043: Data = 4'h2; //+ 
    18'h10044: Data = 4'h2; //+ 
    18'h10045: Data = 4'h2; //+ 
    18'h10046: Data = 4'h2; //+ 
    18'h10047: Data = 4'h2; //+ 
    18'h10048: Data = 4'h2; //+ 
    18'h10049: Data = 4'h4; //> 
    18'h10050: Data = 4'h3; //- 
    18'h10051: Data = 4'h3; //- 
    18'h10052: Data = 4'h3; //- 
    18'h10053: Data = 4'h4; //> 
    18'h10054: Data = 4'h4; //> 
    18'h10055: Data = 4'h4; //> 
    18'h10056: Data = 4'h4; //> 
    18'h10057: Data = 4'h4; //> 
    18'h10058: Data = 4'h4; //> 
    18'h10059: Data = 4'h4; //> 
    18'h10060: Data = 4'h4; //> 
    18'h10061: Data = 4'h4; //> 
    18'h10062: Data = 4'h4; //> 
    18'h10063: Data = 4'h2; //+ 
    18'h10064: Data = 4'h2; //+ 
    18'h10065: Data = 4'h2; //+ 
    18'h10066: Data = 4'h2; //+ 
    18'h10067: Data = 4'h2; //+ 
    18'h10068: Data = 4'h2; //+ 
    18'h10069: Data = 4'h2; //+ 
    18'h10070: Data = 4'h2; //+ 
    18'h10071: Data = 4'h2; //+ 
    18'h10072: Data = 4'h2; //+ 
    18'h10073: Data = 4'h2; //+ 
    18'h10074: Data = 4'h2; //+ 
    18'h10075: Data = 4'h2; //+ 
    18'h10076: Data = 4'h2; //+ 
    18'h10077: Data = 4'h2; //+ 
    18'h10078: Data = 4'h6; //[ 
    18'h10079: Data = 4'h6; //[ 
    18'h10080: Data = 4'h4; //> 
    18'h10081: Data = 4'h4; //> 
    18'h10082: Data = 4'h4; //> 
    18'h10083: Data = 4'h4; //> 
    18'h10084: Data = 4'h4; //> 
    18'h10085: Data = 4'h4; //> 
    18'h10086: Data = 4'h4; //> 
    18'h10087: Data = 4'h4; //> 
    18'h10088: Data = 4'h4; //> 
    18'h10089: Data = 4'h7; //] 
    18'h10090: Data = 4'h2; //+ 
    18'h10091: Data = 4'h6; //[ 
    18'h10092: Data = 4'h5; //< 
    18'h10093: Data = 4'h5; //< 
    18'h10094: Data = 4'h5; //< 
    18'h10095: Data = 4'h5; //< 
    18'h10096: Data = 4'h5; //< 
    18'h10097: Data = 4'h5; //< 
    18'h10098: Data = 4'h5; //< 
    18'h10099: Data = 4'h5; //< 
    18'h10100: Data = 4'h5; //< 
    18'h10101: Data = 4'h7; //] 
    18'h10102: Data = 4'h4; //> 
    18'h10103: Data = 4'h4; //> 
    18'h10104: Data = 4'h4; //> 
    18'h10105: Data = 4'h4; //> 
    18'h10106: Data = 4'h4; //> 
    18'h10107: Data = 4'h4; //> 
    18'h10108: Data = 4'h4; //> 
    18'h10109: Data = 4'h4; //> 
    18'h10110: Data = 4'h4; //> 
    18'h10111: Data = 4'h3; //- 
    18'h10112: Data = 4'h7; //] 
    18'h10113: Data = 4'h2; //+ 
    18'h10114: Data = 4'h6; //[ 
    18'h10115: Data = 4'h4; //> 
    18'h10116: Data = 4'h4; //> 
    18'h10117: Data = 4'h4; //> 
    18'h10118: Data = 4'h4; //> 
    18'h10119: Data = 4'h4; //> 
    18'h10120: Data = 4'h4; //> 
    18'h10121: Data = 4'h4; //> 
    18'h10122: Data = 4'h4; //> 
    18'h10123: Data = 4'ha; //0 
    18'h10124: Data = 4'h4; //> 
    18'h10125: Data = 4'h7; //] 
    18'h10126: Data = 4'h5; //< 
    18'h10127: Data = 4'h5; //< 
    18'h10128: Data = 4'h5; //< 
    18'h10129: Data = 4'h5; //< 
    18'h10130: Data = 4'h5; //< 
    18'h10131: Data = 4'h5; //< 
    18'h10132: Data = 4'h5; //< 
    18'h10133: Data = 4'h5; //< 
    18'h10134: Data = 4'h5; //< 
    18'h10135: Data = 4'h6; //[ 
    18'h10136: Data = 4'h5; //< 
    18'h10137: Data = 4'h5; //< 
    18'h10138: Data = 4'h5; //< 
    18'h10139: Data = 4'h5; //< 
    18'h10140: Data = 4'h5; //< 
    18'h10141: Data = 4'h5; //< 
    18'h10142: Data = 4'h5; //< 
    18'h10143: Data = 4'h5; //< 
    18'h10144: Data = 4'h5; //< 
    18'h10145: Data = 4'h7; //] 
    18'h10146: Data = 4'h4; //> 
    18'h10147: Data = 4'h4; //> 
    18'h10148: Data = 4'h4; //> 
    18'h10149: Data = 4'h4; //> 
    18'h10150: Data = 4'h4; //> 
    18'h10151: Data = 4'h4; //> 
    18'h10152: Data = 4'h4; //> 
    18'h10153: Data = 4'h4; //> 
    18'h10154: Data = 4'ha; //0 
    18'h10155: Data = 4'h2; //+ 
    18'h10156: Data = 4'h5; //< 
    18'h10157: Data = 4'h5; //< 
    18'h10158: Data = 4'h5; //< 
    18'h10159: Data = 4'h5; //< 
    18'h10160: Data = 4'h5; //< 
    18'h10161: Data = 4'h5; //< 
    18'h10162: Data = 4'h5; //< 
    18'h10163: Data = 4'h2; //+ 
    18'h10164: Data = 4'h2; //+ 
    18'h10165: Data = 4'h2; //+ 
    18'h10166: Data = 4'h2; //+ 
    18'h10167: Data = 4'h2; //+ 
    18'h10168: Data = 4'h6; //[ 
    18'h10169: Data = 4'h3; //- 
    18'h10170: Data = 4'h6; //[ 
    18'h10171: Data = 4'h3; //- 
    18'h10172: Data = 4'h4; //> 
    18'h10173: Data = 4'h4; //> 
    18'h10174: Data = 4'h4; //> 
    18'h10175: Data = 4'h4; //> 
    18'h10176: Data = 4'h4; //> 
    18'h10177: Data = 4'h4; //> 
    18'h10178: Data = 4'h4; //> 
    18'h10179: Data = 4'h4; //> 
    18'h10180: Data = 4'h4; //> 
    18'h10181: Data = 4'h2; //+ 
    18'h10182: Data = 4'h5; //< 
    18'h10183: Data = 4'h5; //< 
    18'h10184: Data = 4'h5; //< 
    18'h10185: Data = 4'h5; //< 
    18'h10186: Data = 4'h5; //< 
    18'h10187: Data = 4'h5; //< 
    18'h10188: Data = 4'h5; //< 
    18'h10189: Data = 4'h5; //< 
    18'h10190: Data = 4'h5; //< 
    18'h10191: Data = 4'h7; //] 
    18'h10192: Data = 4'h4; //> 
    18'h10193: Data = 4'h4; //> 
    18'h10194: Data = 4'h4; //> 
    18'h10195: Data = 4'h4; //> 
    18'h10196: Data = 4'h4; //> 
    18'h10197: Data = 4'h4; //> 
    18'h10198: Data = 4'h4; //> 
    18'h10199: Data = 4'h4; //> 
    18'h10200: Data = 4'h4; //> 
    18'h10201: Data = 4'h7; //] 
    18'h10202: Data = 4'h4; //> 
    18'h10203: Data = 4'h4; //> 
    18'h10204: Data = 4'h4; //> 
    18'h10205: Data = 4'h4; //> 
    18'h10206: Data = 4'h4; //> 
    18'h10207: Data = 4'h4; //> 
    18'h10208: Data = 4'h4; //> 
    18'h10209: Data = 4'h2; //+ 
    18'h10210: Data = 4'h4; //> 
    18'h10211: Data = 4'h4; //> 
    18'h10212: Data = 4'h4; //> 
    18'h10213: Data = 4'h4; //> 
    18'h10214: Data = 4'h4; //> 
    18'h10215: Data = 4'h4; //> 
    18'h10216: Data = 4'h4; //> 
    18'h10217: Data = 4'h4; //> 
    18'h10218: Data = 4'h4; //> 
    18'h10219: Data = 4'h4; //> 
    18'h10220: Data = 4'h4; //> 
    18'h10221: Data = 4'h4; //> 
    18'h10222: Data = 4'h4; //> 
    18'h10223: Data = 4'h4; //> 
    18'h10224: Data = 4'h4; //> 
    18'h10225: Data = 4'h4; //> 
    18'h10226: Data = 4'h4; //> 
    18'h10227: Data = 4'h4; //> 
    18'h10228: Data = 4'h4; //> 
    18'h10229: Data = 4'h4; //> 
    18'h10230: Data = 4'h4; //> 
    18'h10231: Data = 4'h4; //> 
    18'h10232: Data = 4'h4; //> 
    18'h10233: Data = 4'h4; //> 
    18'h10234: Data = 4'h4; //> 
    18'h10235: Data = 4'h4; //> 
    18'h10236: Data = 4'h4; //> 
    18'h10237: Data = 4'h2; //+ 
    18'h10238: Data = 4'h5; //< 
    18'h10239: Data = 4'h5; //< 
    18'h10240: Data = 4'h5; //< 
    18'h10241: Data = 4'h5; //< 
    18'h10242: Data = 4'h5; //< 
    18'h10243: Data = 4'h5; //< 
    18'h10244: Data = 4'h5; //< 
    18'h10245: Data = 4'h5; //< 
    18'h10246: Data = 4'h5; //< 
    18'h10247: Data = 4'h5; //< 
    18'h10248: Data = 4'h5; //< 
    18'h10249: Data = 4'h5; //< 
    18'h10250: Data = 4'h5; //< 
    18'h10251: Data = 4'h5; //< 
    18'h10252: Data = 4'h5; //< 
    18'h10253: Data = 4'h5; //< 
    18'h10254: Data = 4'h5; //< 
    18'h10255: Data = 4'h6; //[ 
    18'h10256: Data = 4'h5; //< 
    18'h10257: Data = 4'h5; //< 
    18'h10258: Data = 4'h5; //< 
    18'h10259: Data = 4'h5; //< 
    18'h10260: Data = 4'h5; //< 
    18'h10261: Data = 4'h5; //< 
    18'h10262: Data = 4'h5; //< 
    18'h10263: Data = 4'h5; //< 
    18'h10264: Data = 4'h5; //< 
    18'h10265: Data = 4'h7; //] 
    18'h10266: Data = 4'h4; //> 
    18'h10267: Data = 4'h4; //> 
    18'h10268: Data = 4'h4; //> 
    18'h10269: Data = 4'ha; //0 
    18'h10270: Data = 4'h2; //+ 
    18'h10271: Data = 4'h6; //[ 
    18'h10272: Data = 4'h4; //> 
    18'h10273: Data = 4'h4; //> 
    18'h10274: Data = 4'h4; //> 
    18'h10275: Data = 4'h4; //> 
    18'h10276: Data = 4'h4; //> 
    18'h10277: Data = 4'h4; //> 
    18'h10278: Data = 4'h6; //[ 
    18'h10279: Data = 4'h4; //> 
    18'h10280: Data = 4'h4; //> 
    18'h10281: Data = 4'h4; //> 
    18'h10282: Data = 4'h4; //> 
    18'h10283: Data = 4'h4; //> 
    18'h10284: Data = 4'h4; //> 
    18'h10285: Data = 4'h4; //> 
    18'h10286: Data = 4'ha; //0 
    18'h10287: Data = 4'h4; //> 
    18'h10288: Data = 4'h4; //> 
    18'h10289: Data = 4'h7; //] 
    18'h10290: Data = 4'h5; //< 
    18'h10291: Data = 4'h5; //< 
    18'h10292: Data = 4'h5; //< 
    18'h10293: Data = 4'h5; //< 
    18'h10294: Data = 4'h5; //< 
    18'h10295: Data = 4'h5; //< 
    18'h10296: Data = 4'h5; //< 
    18'h10297: Data = 4'h5; //< 
    18'h10298: Data = 4'h5; //< 
    18'h10299: Data = 4'h6; //[ 
    18'h10300: Data = 4'h5; //< 
    18'h10301: Data = 4'h5; //< 
    18'h10302: Data = 4'h5; //< 
    18'h10303: Data = 4'h5; //< 
    18'h10304: Data = 4'h5; //< 
    18'h10305: Data = 4'h5; //< 
    18'h10306: Data = 4'h5; //< 
    18'h10307: Data = 4'h5; //< 
    18'h10308: Data = 4'h5; //< 
    18'h10309: Data = 4'h7; //] 
    18'h10310: Data = 4'h4; //> 
    18'h10311: Data = 4'h4; //> 
    18'h10312: Data = 4'h4; //> 
    18'h10313: Data = 4'h4; //> 
    18'h10314: Data = 4'h4; //> 
    18'h10315: Data = 4'h4; //> 
    18'h10316: Data = 4'h4; //> 
    18'h10317: Data = 4'ha; //0 
    18'h10318: Data = 4'h2; //+ 
    18'h10319: Data = 4'h5; //< 
    18'h10320: Data = 4'h5; //< 
    18'h10321: Data = 4'h5; //< 
    18'h10322: Data = 4'h5; //< 
    18'h10323: Data = 4'h5; //< 
    18'h10324: Data = 4'h5; //< 
    18'h10325: Data = 4'h2; //+ 
    18'h10326: Data = 4'h2; //+ 
    18'h10327: Data = 4'h2; //+ 
    18'h10328: Data = 4'h2; //+ 
    18'h10329: Data = 4'h6; //[ 
    18'h10330: Data = 4'h3; //- 
    18'h10331: Data = 4'h6; //[ 
    18'h10332: Data = 4'h3; //- 
    18'h10333: Data = 4'h4; //> 
    18'h10334: Data = 4'h4; //> 
    18'h10335: Data = 4'h4; //> 
    18'h10336: Data = 4'h4; //> 
    18'h10337: Data = 4'h4; //> 
    18'h10338: Data = 4'h4; //> 
    18'h10339: Data = 4'h4; //> 
    18'h10340: Data = 4'h4; //> 
    18'h10341: Data = 4'h4; //> 
    18'h10342: Data = 4'h2; //+ 
    18'h10343: Data = 4'h5; //< 
    18'h10344: Data = 4'h5; //< 
    18'h10345: Data = 4'h5; //< 
    18'h10346: Data = 4'h5; //< 
    18'h10347: Data = 4'h5; //< 
    18'h10348: Data = 4'h5; //< 
    18'h10349: Data = 4'h5; //< 
    18'h10350: Data = 4'h5; //< 
    18'h10351: Data = 4'h5; //< 
    18'h10352: Data = 4'h7; //] 
    18'h10353: Data = 4'h4; //> 
    18'h10354: Data = 4'h4; //> 
    18'h10355: Data = 4'h4; //> 
    18'h10356: Data = 4'h4; //> 
    18'h10357: Data = 4'h4; //> 
    18'h10358: Data = 4'h4; //> 
    18'h10359: Data = 4'h4; //> 
    18'h10360: Data = 4'h4; //> 
    18'h10361: Data = 4'h4; //> 
    18'h10362: Data = 4'h7; //] 
    18'h10363: Data = 4'h4; //> 
    18'h10364: Data = 4'h4; //> 
    18'h10365: Data = 4'h4; //> 
    18'h10366: Data = 4'h4; //> 
    18'h10367: Data = 4'h4; //> 
    18'h10368: Data = 4'h4; //> 
    18'h10369: Data = 4'h2; //+ 
    18'h10370: Data = 4'h5; //< 
    18'h10371: Data = 4'h5; //< 
    18'h10372: Data = 4'h5; //< 
    18'h10373: Data = 4'h5; //< 
    18'h10374: Data = 4'h5; //< 
    18'h10375: Data = 4'h5; //< 
    18'h10376: Data = 4'h2; //+ 
    18'h10377: Data = 4'h2; //+ 
    18'h10378: Data = 4'h2; //+ 
    18'h10379: Data = 4'h2; //+ 
    18'h10380: Data = 4'h2; //+ 
    18'h10381: Data = 4'h2; //+ 
    18'h10382: Data = 4'h2; //+ 
    18'h10383: Data = 4'h6; //[ 
    18'h10384: Data = 4'h3; //- 
    18'h10385: Data = 4'h6; //[ 
    18'h10386: Data = 4'h3; //- 
    18'h10387: Data = 4'h4; //> 
    18'h10388: Data = 4'h4; //> 
    18'h10389: Data = 4'h4; //> 
    18'h10390: Data = 4'h4; //> 
    18'h10391: Data = 4'h4; //> 
    18'h10392: Data = 4'h4; //> 
    18'h10393: Data = 4'h4; //> 
    18'h10394: Data = 4'h4; //> 
    18'h10395: Data = 4'h4; //> 
    18'h10396: Data = 4'h2; //+ 
    18'h10397: Data = 4'h5; //< 
    18'h10398: Data = 4'h5; //< 
    18'h10399: Data = 4'h5; //< 
    18'h10400: Data = 4'h5; //< 
    18'h10401: Data = 4'h5; //< 
    18'h10402: Data = 4'h5; //< 
    18'h10403: Data = 4'h5; //< 
    18'h10404: Data = 4'h5; //< 
    18'h10405: Data = 4'h5; //< 
    18'h10406: Data = 4'h7; //] 
    18'h10407: Data = 4'h4; //> 
    18'h10408: Data = 4'h4; //> 
    18'h10409: Data = 4'h4; //> 
    18'h10410: Data = 4'h4; //> 
    18'h10411: Data = 4'h4; //> 
    18'h10412: Data = 4'h4; //> 
    18'h10413: Data = 4'h4; //> 
    18'h10414: Data = 4'h4; //> 
    18'h10415: Data = 4'h4; //> 
    18'h10416: Data = 4'h7; //] 
    18'h10417: Data = 4'h4; //> 
    18'h10418: Data = 4'h4; //> 
    18'h10419: Data = 4'h4; //> 
    18'h10420: Data = 4'h4; //> 
    18'h10421: Data = 4'h4; //> 
    18'h10422: Data = 4'h4; //> 
    18'h10423: Data = 4'h2; //+ 
    18'h10424: Data = 4'h5; //< 
    18'h10425: Data = 4'h5; //< 
    18'h10426: Data = 4'h5; //< 
    18'h10427: Data = 4'h5; //< 
    18'h10428: Data = 4'h5; //< 
    18'h10429: Data = 4'h5; //< 
    18'h10430: Data = 4'h5; //< 
    18'h10431: Data = 4'h5; //< 
    18'h10432: Data = 4'h5; //< 
    18'h10433: Data = 4'h5; //< 
    18'h10434: Data = 4'h5; //< 
    18'h10435: Data = 4'h5; //< 
    18'h10436: Data = 4'h5; //< 
    18'h10437: Data = 4'h5; //< 
    18'h10438: Data = 4'h5; //< 
    18'h10439: Data = 4'h5; //< 
    18'h10440: Data = 4'h6; //[ 
    18'h10441: Data = 4'h5; //< 
    18'h10442: Data = 4'h5; //< 
    18'h10443: Data = 4'h5; //< 
    18'h10444: Data = 4'h5; //< 
    18'h10445: Data = 4'h5; //< 
    18'h10446: Data = 4'h5; //< 
    18'h10447: Data = 4'h5; //< 
    18'h10448: Data = 4'h5; //< 
    18'h10449: Data = 4'h5; //< 
    18'h10450: Data = 4'h7; //] 
    18'h10451: Data = 4'h4; //> 
    18'h10452: Data = 4'h4; //> 
    18'h10453: Data = 4'h4; //> 
    18'h10454: Data = 4'h6; //[ 
    18'h10455: Data = 4'ha; //0 
    18'h10456: Data = 4'h4; //> 
    18'h10457: Data = 4'h4; //> 
    18'h10458: Data = 4'h4; //> 
    18'h10459: Data = 4'h4; //> 
    18'h10460: Data = 4'h4; //> 
    18'h10461: Data = 4'h4; //> 
    18'h10462: Data = 4'h6; //[ 
    18'h10463: Data = 4'h4; //> 
    18'h10464: Data = 4'h4; //> 
    18'h10465: Data = 4'h4; //> 
    18'h10466: Data = 4'h4; //> 
    18'h10467: Data = 4'h4; //> 
    18'h10468: Data = 4'h4; //> 
    18'h10469: Data = 4'h4; //> 
    18'h10470: Data = 4'h6; //[ 
    18'h10471: Data = 4'h3; //- 
    18'h10472: Data = 4'h5; //< 
    18'h10473: Data = 4'h5; //< 
    18'h10474: Data = 4'h5; //< 
    18'h10475: Data = 4'h5; //< 
    18'h10476: Data = 4'h5; //< 
    18'h10477: Data = 4'h5; //< 
    18'h10478: Data = 4'h2; //+ 
    18'h10479: Data = 4'h4; //> 
    18'h10480: Data = 4'h4; //> 
    18'h10481: Data = 4'h4; //> 
    18'h10482: Data = 4'h4; //> 
    18'h10483: Data = 4'h4; //> 
    18'h10484: Data = 4'h4; //> 
    18'h10485: Data = 4'h7; //] 
    18'h10486: Data = 4'h5; //< 
    18'h10487: Data = 4'h5; //< 
    18'h10488: Data = 4'h5; //< 
    18'h10489: Data = 4'h5; //< 
    18'h10490: Data = 4'h5; //< 
    18'h10491: Data = 4'h5; //< 
    18'h10492: Data = 4'h6; //[ 
    18'h10493: Data = 4'h3; //- 
    18'h10494: Data = 4'h4; //> 
    18'h10495: Data = 4'h4; //> 
    18'h10496: Data = 4'h4; //> 
    18'h10497: Data = 4'h4; //> 
    18'h10498: Data = 4'h4; //> 
    18'h10499: Data = 4'h4; //> 
    18'h10500: Data = 4'h2; //+ 
    18'h10501: Data = 4'h5; //< 
    18'h10502: Data = 4'h5; //< 
    18'h10503: Data = 4'h2; //+ 
    18'h10504: Data = 4'h5; //< 
    18'h10505: Data = 4'h5; //< 
    18'h10506: Data = 4'h5; //< 
    18'h10507: Data = 4'h2; //+ 
    18'h10508: Data = 4'h5; //< 
    18'h10509: Data = 4'h7; //] 
    18'h10510: Data = 4'h4; //> 
    18'h10511: Data = 4'h4; //> 
    18'h10512: Data = 4'h4; //> 
    18'h10513: Data = 4'h4; //> 
    18'h10514: Data = 4'h4; //> 
    18'h10515: Data = 4'h4; //> 
    18'h10516: Data = 4'h4; //> 
    18'h10517: Data = 4'h4; //> 
    18'h10518: Data = 4'h7; //] 
    18'h10519: Data = 4'h5; //< 
    18'h10520: Data = 4'h5; //< 
    18'h10521: Data = 4'h5; //< 
    18'h10522: Data = 4'h5; //< 
    18'h10523: Data = 4'h5; //< 
    18'h10524: Data = 4'h5; //< 
    18'h10525: Data = 4'h5; //< 
    18'h10526: Data = 4'h5; //< 
    18'h10527: Data = 4'h5; //< 
    18'h10528: Data = 4'h6; //[ 
    18'h10529: Data = 4'h5; //< 
    18'h10530: Data = 4'h5; //< 
    18'h10531: Data = 4'h5; //< 
    18'h10532: Data = 4'h5; //< 
    18'h10533: Data = 4'h5; //< 
    18'h10534: Data = 4'h5; //< 
    18'h10535: Data = 4'h5; //< 
    18'h10536: Data = 4'h5; //< 
    18'h10537: Data = 4'h5; //< 
    18'h10538: Data = 4'h7; //] 
    18'h10539: Data = 4'h4; //> 
    18'h10540: Data = 4'h4; //> 
    18'h10541: Data = 4'h4; //> 
    18'h10542: Data = 4'h4; //> 
    18'h10543: Data = 4'h4; //> 
    18'h10544: Data = 4'h4; //> 
    18'h10545: Data = 4'h4; //> 
    18'h10546: Data = 4'h4; //> 
    18'h10547: Data = 4'h4; //> 
    18'h10548: Data = 4'h6; //[ 
    18'h10549: Data = 4'h4; //> 
    18'h10550: Data = 4'h4; //> 
    18'h10551: Data = 4'h4; //> 
    18'h10552: Data = 4'h4; //> 
    18'h10553: Data = 4'h4; //> 
    18'h10554: Data = 4'h4; //> 
    18'h10555: Data = 4'h4; //> 
    18'h10556: Data = 4'h4; //> 
    18'h10557: Data = 4'h6; //[ 
    18'h10558: Data = 4'h3; //- 
    18'h10559: Data = 4'h5; //< 
    18'h10560: Data = 4'h5; //< 
    18'h10561: Data = 4'h5; //< 
    18'h10562: Data = 4'h5; //< 
    18'h10563: Data = 4'h5; //< 
    18'h10564: Data = 4'h5; //< 
    18'h10565: Data = 4'h5; //< 
    18'h10566: Data = 4'h2; //+ 
    18'h10567: Data = 4'h4; //> 
    18'h10568: Data = 4'h4; //> 
    18'h10569: Data = 4'h4; //> 
    18'h10570: Data = 4'h4; //> 
    18'h10571: Data = 4'h4; //> 
    18'h10572: Data = 4'h4; //> 
    18'h10573: Data = 4'h4; //> 
    18'h10574: Data = 4'h7; //] 
    18'h10575: Data = 4'h5; //< 
    18'h10576: Data = 4'h5; //< 
    18'h10577: Data = 4'h5; //< 
    18'h10578: Data = 4'h5; //< 
    18'h10579: Data = 4'h5; //< 
    18'h10580: Data = 4'h5; //< 
    18'h10581: Data = 4'h5; //< 
    18'h10582: Data = 4'h6; //[ 
    18'h10583: Data = 4'h3; //- 
    18'h10584: Data = 4'h4; //> 
    18'h10585: Data = 4'h4; //> 
    18'h10586: Data = 4'h4; //> 
    18'h10587: Data = 4'h4; //> 
    18'h10588: Data = 4'h4; //> 
    18'h10589: Data = 4'h4; //> 
    18'h10590: Data = 4'h4; //> 
    18'h10591: Data = 4'h2; //+ 
    18'h10592: Data = 4'h5; //< 
    18'h10593: Data = 4'h5; //< 
    18'h10594: Data = 4'h2; //+ 
    18'h10595: Data = 4'h5; //< 
    18'h10596: Data = 4'h5; //< 
    18'h10597: Data = 4'h5; //< 
    18'h10598: Data = 4'h2; //+ 
    18'h10599: Data = 4'h5; //< 
    18'h10600: Data = 4'h5; //< 
    18'h10601: Data = 4'h7; //] 
    18'h10602: Data = 4'h4; //> 
    18'h10603: Data = 4'h4; //> 
    18'h10604: Data = 4'h4; //> 
    18'h10605: Data = 4'h4; //> 
    18'h10606: Data = 4'h4; //> 
    18'h10607: Data = 4'h4; //> 
    18'h10608: Data = 4'h4; //> 
    18'h10609: Data = 4'h4; //> 
    18'h10610: Data = 4'h7; //] 
    18'h10611: Data = 4'h5; //< 
    18'h10612: Data = 4'h5; //< 
    18'h10613: Data = 4'h5; //< 
    18'h10614: Data = 4'h5; //< 
    18'h10615: Data = 4'h5; //< 
    18'h10616: Data = 4'h5; //< 
    18'h10617: Data = 4'h5; //< 
    18'h10618: Data = 4'h5; //< 
    18'h10619: Data = 4'h5; //< 
    18'h10620: Data = 4'h6; //[ 
    18'h10621: Data = 4'h5; //< 
    18'h10622: Data = 4'h5; //< 
    18'h10623: Data = 4'h5; //< 
    18'h10624: Data = 4'h5; //< 
    18'h10625: Data = 4'h5; //< 
    18'h10626: Data = 4'h5; //< 
    18'h10627: Data = 4'h5; //< 
    18'h10628: Data = 4'h5; //< 
    18'h10629: Data = 4'h5; //< 
    18'h10630: Data = 4'h7; //] 
    18'h10631: Data = 4'h4; //> 
    18'h10632: Data = 4'h4; //> 
    18'h10633: Data = 4'h4; //> 
    18'h10634: Data = 4'h4; //> 
    18'h10635: Data = 4'h4; //> 
    18'h10636: Data = 4'h4; //> 
    18'h10637: Data = 4'h4; //> 
    18'h10638: Data = 4'h6; //[ 
    18'h10639: Data = 4'h3; //- 
    18'h10640: Data = 4'h5; //< 
    18'h10641: Data = 4'h5; //< 
    18'h10642: Data = 4'h5; //< 
    18'h10643: Data = 4'h5; //< 
    18'h10644: Data = 4'h5; //< 
    18'h10645: Data = 4'h5; //< 
    18'h10646: Data = 4'h5; //< 
    18'h10647: Data = 4'h2; //+ 
    18'h10648: Data = 4'h4; //> 
    18'h10649: Data = 4'h4; //> 
    18'h10650: Data = 4'h4; //> 
    18'h10651: Data = 4'h4; //> 
    18'h10652: Data = 4'h4; //> 
    18'h10653: Data = 4'h4; //> 
    18'h10654: Data = 4'h4; //> 
    18'h10655: Data = 4'h7; //] 
    18'h10656: Data = 4'h5; //< 
    18'h10657: Data = 4'h5; //< 
    18'h10658: Data = 4'h5; //< 
    18'h10659: Data = 4'h5; //< 
    18'h10660: Data = 4'h5; //< 
    18'h10661: Data = 4'h5; //< 
    18'h10662: Data = 4'h5; //< 
    18'h10663: Data = 4'h6; //[ 
    18'h10664: Data = 4'h3; //- 
    18'h10665: Data = 4'h4; //> 
    18'h10666: Data = 4'h4; //> 
    18'h10667: Data = 4'h4; //> 
    18'h10668: Data = 4'h4; //> 
    18'h10669: Data = 4'h4; //> 
    18'h10670: Data = 4'h4; //> 
    18'h10671: Data = 4'h4; //> 
    18'h10672: Data = 4'h2; //+ 
    18'h10673: Data = 4'h5; //< 
    18'h10674: Data = 4'h5; //< 
    18'h10675: Data = 4'h2; //+ 
    18'h10676: Data = 4'h5; //< 
    18'h10677: Data = 4'h5; //< 
    18'h10678: Data = 4'h5; //< 
    18'h10679: Data = 4'h5; //< 
    18'h10680: Data = 4'h5; //< 
    18'h10681: Data = 4'h7; //] 
    18'h10682: Data = 4'h4; //> 
    18'h10683: Data = 4'h4; //> 
    18'h10684: Data = 4'h4; //> 
    18'h10685: Data = 4'h4; //> 
    18'h10686: Data = 4'h4; //> 
    18'h10687: Data = 4'h4; //> 
    18'h10688: Data = 4'h4; //> 
    18'h10689: Data = 4'h4; //> 
    18'h10690: Data = 4'h4; //> 
    18'h10691: Data = 4'h2; //+ 
    18'h10692: Data = 4'h2; //+ 
    18'h10693: Data = 4'h2; //+ 
    18'h10694: Data = 4'h2; //+ 
    18'h10695: Data = 4'h2; //+ 
    18'h10696: Data = 4'h2; //+ 
    18'h10697: Data = 4'h2; //+ 
    18'h10698: Data = 4'h2; //+ 
    18'h10699: Data = 4'h2; //+ 
    18'h10700: Data = 4'h2; //+ 
    18'h10701: Data = 4'h2; //+ 
    18'h10702: Data = 4'h2; //+ 
    18'h10703: Data = 4'h2; //+ 
    18'h10704: Data = 4'h2; //+ 
    18'h10705: Data = 4'h2; //+ 
    18'h10706: Data = 4'h6; //[ 
    18'h10707: Data = 4'h6; //[ 
    18'h10708: Data = 4'h4; //> 
    18'h10709: Data = 4'h4; //> 
    18'h10710: Data = 4'h4; //> 
    18'h10711: Data = 4'h4; //> 
    18'h10712: Data = 4'h4; //> 
    18'h10713: Data = 4'h4; //> 
    18'h10714: Data = 4'h4; //> 
    18'h10715: Data = 4'h4; //> 
    18'h10716: Data = 4'h4; //> 
    18'h10717: Data = 4'h7; //] 
    18'h10718: Data = 4'h2; //+ 
    18'h10719: Data = 4'h4; //> 
    18'h10720: Data = 4'ha; //0 
    18'h10721: Data = 4'h4; //> 
    18'h10722: Data = 4'ha; //0 
    18'h10723: Data = 4'h4; //> 
    18'h10724: Data = 4'ha; //0 
    18'h10725: Data = 4'h4; //> 
    18'h10726: Data = 4'ha; //0 
    18'h10727: Data = 4'h4; //> 
    18'h10728: Data = 4'ha; //0 
    18'h10729: Data = 4'h4; //> 
    18'h10730: Data = 4'ha; //0 
    18'h10731: Data = 4'h4; //> 
    18'h10732: Data = 4'ha; //0 
    18'h10733: Data = 4'h4; //> 
    18'h10734: Data = 4'ha; //0 
    18'h10735: Data = 4'h4; //> 
    18'h10736: Data = 4'ha; //0 
    18'h10737: Data = 4'h5; //< 
    18'h10738: Data = 4'h5; //< 
    18'h10739: Data = 4'h5; //< 
    18'h10740: Data = 4'h5; //< 
    18'h10741: Data = 4'h5; //< 
    18'h10742: Data = 4'h5; //< 
    18'h10743: Data = 4'h5; //< 
    18'h10744: Data = 4'h5; //< 
    18'h10745: Data = 4'h5; //< 
    18'h10746: Data = 4'h6; //[ 
    18'h10747: Data = 4'h5; //< 
    18'h10748: Data = 4'h5; //< 
    18'h10749: Data = 4'h5; //< 
    18'h10750: Data = 4'h5; //< 
    18'h10751: Data = 4'h5; //< 
    18'h10752: Data = 4'h5; //< 
    18'h10753: Data = 4'h5; //< 
    18'h10754: Data = 4'h5; //< 
    18'h10755: Data = 4'h5; //< 
    18'h10756: Data = 4'h7; //] 
    18'h10757: Data = 4'h4; //> 
    18'h10758: Data = 4'h4; //> 
    18'h10759: Data = 4'h4; //> 
    18'h10760: Data = 4'h4; //> 
    18'h10761: Data = 4'h4; //> 
    18'h10762: Data = 4'h4; //> 
    18'h10763: Data = 4'h4; //> 
    18'h10764: Data = 4'h4; //> 
    18'h10765: Data = 4'h4; //> 
    18'h10766: Data = 4'h3; //- 
    18'h10767: Data = 4'h7; //] 
    18'h10768: Data = 4'h2; //+ 
    18'h10769: Data = 4'h6; //[ 
    18'h10770: Data = 4'h4; //> 
    18'h10771: Data = 4'h2; //+ 
    18'h10772: Data = 4'h4; //> 
    18'h10773: Data = 4'h4; //> 
    18'h10774: Data = 4'h4; //> 
    18'h10775: Data = 4'h4; //> 
    18'h10776: Data = 4'h4; //> 
    18'h10777: Data = 4'h4; //> 
    18'h10778: Data = 4'h4; //> 
    18'h10779: Data = 4'h4; //> 
    18'h10780: Data = 4'h7; //] 
    18'h10781: Data = 4'h5; //< 
    18'h10782: Data = 4'h5; //< 
    18'h10783: Data = 4'h5; //< 
    18'h10784: Data = 4'h5; //< 
    18'h10785: Data = 4'h5; //< 
    18'h10786: Data = 4'h5; //< 
    18'h10787: Data = 4'h5; //< 
    18'h10788: Data = 4'h5; //< 
    18'h10789: Data = 4'h5; //< 
    18'h10790: Data = 4'h6; //[ 
    18'h10791: Data = 4'h5; //< 
    18'h10792: Data = 4'h5; //< 
    18'h10793: Data = 4'h5; //< 
    18'h10794: Data = 4'h5; //< 
    18'h10795: Data = 4'h5; //< 
    18'h10796: Data = 4'h5; //< 
    18'h10797: Data = 4'h5; //< 
    18'h10798: Data = 4'h5; //< 
    18'h10799: Data = 4'h5; //< 
    18'h10800: Data = 4'h7; //] 
    18'h10801: Data = 4'h4; //> 
    18'h10802: Data = 4'h4; //> 
    18'h10803: Data = 4'h4; //> 
    18'h10804: Data = 4'h4; //> 
    18'h10805: Data = 4'h4; //> 
    18'h10806: Data = 4'h4; //> 
    18'h10807: Data = 4'h4; //> 
    18'h10808: Data = 4'h4; //> 
    18'h10809: Data = 4'h4; //> 
    18'h10810: Data = 4'h6; //[ 
    18'h10811: Data = 4'h4; //> 
    18'h10812: Data = 4'h3; //- 
    18'h10813: Data = 4'h4; //> 
    18'h10814: Data = 4'h4; //> 
    18'h10815: Data = 4'h4; //> 
    18'h10816: Data = 4'h4; //> 
    18'h10817: Data = 4'h6; //[ 
    18'h10818: Data = 4'h3; //- 
    18'h10819: Data = 4'h5; //< 
    18'h10820: Data = 4'h5; //< 
    18'h10821: Data = 4'h5; //< 
    18'h10822: Data = 4'h5; //< 
    18'h10823: Data = 4'h2; //+ 
    18'h10824: Data = 4'h4; //> 
    18'h10825: Data = 4'h4; //> 
    18'h10826: Data = 4'h4; //> 
    18'h10827: Data = 4'h4; //> 
    18'h10828: Data = 4'h7; //] 
    18'h10829: Data = 4'h5; //< 
    18'h10830: Data = 4'h5; //< 
    18'h10831: Data = 4'h5; //< 
    18'h10832: Data = 4'h5; //< 
    18'h10833: Data = 4'h6; //[ 
    18'h10834: Data = 4'h3; //- 
    18'h10835: Data = 4'h4; //> 
    18'h10836: Data = 4'h4; //> 
    18'h10837: Data = 4'h4; //> 
    18'h10838: Data = 4'h4; //> 
    18'h10839: Data = 4'h2; //+ 
    18'h10840: Data = 4'h5; //< 
    18'h10841: Data = 4'h5; //< 
    18'h10842: Data = 4'h5; //< 
    18'h10843: Data = 4'h5; //< 
    18'h10844: Data = 4'h5; //< 
    18'h10845: Data = 4'h6; //[ 
    18'h10846: Data = 4'h3; //- 
    18'h10847: Data = 4'h4; //> 
    18'h10848: Data = 4'h4; //> 
    18'h10849: Data = 4'h6; //[ 
    18'h10850: Data = 4'h3; //- 
    18'h10851: Data = 4'h5; //< 
    18'h10852: Data = 4'h5; //< 
    18'h10853: Data = 4'h2; //+ 
    18'h10854: Data = 4'h4; //> 
    18'h10855: Data = 4'h4; //> 
    18'h10856: Data = 4'h7; //] 
    18'h10857: Data = 4'h5; //< 
    18'h10858: Data = 4'h5; //< 
    18'h10859: Data = 4'h6; //[ 
    18'h10860: Data = 4'h3; //- 
    18'h10861: Data = 4'h4; //> 
    18'h10862: Data = 4'h4; //> 
    18'h10863: Data = 4'h2; //+ 
    18'h10864: Data = 4'h4; //> 
    18'h10865: Data = 4'h4; //> 
    18'h10866: Data = 4'h2; //+ 
    18'h10867: Data = 4'h5; //< 
    18'h10868: Data = 4'h5; //< 
    18'h10869: Data = 4'h5; //< 
    18'h10870: Data = 4'h5; //< 
    18'h10871: Data = 4'h7; //] 
    18'h10872: Data = 4'h2; //+ 
    18'h10873: Data = 4'h4; //> 
    18'h10874: Data = 4'h4; //> 
    18'h10875: Data = 4'h4; //> 
    18'h10876: Data = 4'h4; //> 
    18'h10877: Data = 4'h4; //> 
    18'h10878: Data = 4'h4; //> 
    18'h10879: Data = 4'h4; //> 
    18'h10880: Data = 4'h4; //> 
    18'h10881: Data = 4'h4; //> 
    18'h10882: Data = 4'h7; //] 
    18'h10883: Data = 4'h5; //< 
    18'h10884: Data = 4'h5; //< 
    18'h10885: Data = 4'h5; //< 
    18'h10886: Data = 4'h5; //< 
    18'h10887: Data = 4'h5; //< 
    18'h10888: Data = 4'h5; //< 
    18'h10889: Data = 4'h5; //< 
    18'h10890: Data = 4'h5; //< 
    18'h10891: Data = 4'h6; //[ 
    18'h10892: Data = 4'h5; //< 
    18'h10893: Data = 4'h5; //< 
    18'h10894: Data = 4'h5; //< 
    18'h10895: Data = 4'h5; //< 
    18'h10896: Data = 4'h5; //< 
    18'h10897: Data = 4'h5; //< 
    18'h10898: Data = 4'h5; //< 
    18'h10899: Data = 4'h5; //< 
    18'h10900: Data = 4'h5; //< 
    18'h10901: Data = 4'h7; //] 
    18'h10902: Data = 4'h7; //] 
    18'h10903: Data = 4'h4; //> 
    18'h10904: Data = 4'h4; //> 
    18'h10905: Data = 4'h4; //> 
    18'h10906: Data = 4'h4; //> 
    18'h10907: Data = 4'h4; //> 
    18'h10908: Data = 4'h4; //> 
    18'h10909: Data = 4'h4; //> 
    18'h10910: Data = 4'h4; //> 
    18'h10911: Data = 4'h4; //> 
    18'h10912: Data = 4'h6; //[ 
    18'h10913: Data = 4'h4; //> 
    18'h10914: Data = 4'h4; //> 
    18'h10915: Data = 4'h4; //> 
    18'h10916: Data = 4'h4; //> 
    18'h10917: Data = 4'h4; //> 
    18'h10918: Data = 4'h4; //> 
    18'h10919: Data = 4'h4; //> 
    18'h10920: Data = 4'h4; //> 
    18'h10921: Data = 4'h4; //> 
    18'h10922: Data = 4'h7; //] 
    18'h10923: Data = 4'h5; //< 
    18'h10924: Data = 4'h5; //< 
    18'h10925: Data = 4'h5; //< 
    18'h10926: Data = 4'h5; //< 
    18'h10927: Data = 4'h5; //< 
    18'h10928: Data = 4'h5; //< 
    18'h10929: Data = 4'h5; //< 
    18'h10930: Data = 4'h5; //< 
    18'h10931: Data = 4'h5; //< 
    18'h10932: Data = 4'h6; //[ 
    18'h10933: Data = 4'h4; //> 
    18'h10934: Data = 4'h6; //[ 
    18'h10935: Data = 4'h3; //- 
    18'h10936: Data = 4'h4; //> 
    18'h10937: Data = 4'h4; //> 
    18'h10938: Data = 4'h4; //> 
    18'h10939: Data = 4'h4; //> 
    18'h10940: Data = 4'h4; //> 
    18'h10941: Data = 4'h4; //> 
    18'h10942: Data = 4'h4; //> 
    18'h10943: Data = 4'h4; //> 
    18'h10944: Data = 4'h4; //> 
    18'h10945: Data = 4'h2; //+ 
    18'h10946: Data = 4'h5; //< 
    18'h10947: Data = 4'h5; //< 
    18'h10948: Data = 4'h5; //< 
    18'h10949: Data = 4'h5; //< 
    18'h10950: Data = 4'h5; //< 
    18'h10951: Data = 4'h5; //< 
    18'h10952: Data = 4'h5; //< 
    18'h10953: Data = 4'h5; //< 
    18'h10954: Data = 4'h5; //< 
    18'h10955: Data = 4'h7; //] 
    18'h10956: Data = 4'h5; //< 
    18'h10957: Data = 4'h5; //< 
    18'h10958: Data = 4'h5; //< 
    18'h10959: Data = 4'h5; //< 
    18'h10960: Data = 4'h5; //< 
    18'h10961: Data = 4'h5; //< 
    18'h10962: Data = 4'h5; //< 
    18'h10963: Data = 4'h5; //< 
    18'h10964: Data = 4'h5; //< 
    18'h10965: Data = 4'h5; //< 
    18'h10966: Data = 4'h7; //] 
    18'h10967: Data = 4'h4; //> 
    18'h10968: Data = 4'h6; //[ 
    18'h10969: Data = 4'h3; //- 
    18'h10970: Data = 4'h4; //> 
    18'h10971: Data = 4'h4; //> 
    18'h10972: Data = 4'h4; //> 
    18'h10973: Data = 4'h4; //> 
    18'h10974: Data = 4'h4; //> 
    18'h10975: Data = 4'h4; //> 
    18'h10976: Data = 4'h4; //> 
    18'h10977: Data = 4'h4; //> 
    18'h10978: Data = 4'h4; //> 
    18'h10979: Data = 4'h2; //+ 
    18'h10980: Data = 4'h5; //< 
    18'h10981: Data = 4'h5; //< 
    18'h10982: Data = 4'h5; //< 
    18'h10983: Data = 4'h5; //< 
    18'h10984: Data = 4'h5; //< 
    18'h10985: Data = 4'h5; //< 
    18'h10986: Data = 4'h5; //< 
    18'h10987: Data = 4'h5; //< 
    18'h10988: Data = 4'h5; //< 
    18'h10989: Data = 4'h7; //] 
    18'h10990: Data = 4'h5; //< 
    18'h10991: Data = 4'h2; //+ 
    18'h10992: Data = 4'h4; //> 
    18'h10993: Data = 4'h4; //> 
    18'h10994: Data = 4'h4; //> 
    18'h10995: Data = 4'h4; //> 
    18'h10996: Data = 4'h4; //> 
    18'h10997: Data = 4'h4; //> 
    18'h10998: Data = 4'h4; //> 
    18'h10999: Data = 4'h4; //> 
    18'h11000: Data = 4'h7; //] 
    18'h11001: Data = 4'h5; //< 
    18'h11002: Data = 4'h5; //< 
    18'h11003: Data = 4'h5; //< 
    18'h11004: Data = 4'h5; //< 
    18'h11005: Data = 4'h5; //< 
    18'h11006: Data = 4'h5; //< 
    18'h11007: Data = 4'h5; //< 
    18'h11008: Data = 4'h5; //< 
    18'h11009: Data = 4'h5; //< 
    18'h11010: Data = 4'h6; //[ 
    18'h11011: Data = 4'h4; //> 
    18'h11012: Data = 4'ha; //0 
    18'h11013: Data = 4'h5; //< 
    18'h11014: Data = 4'h3; //- 
    18'h11015: Data = 4'h4; //> 
    18'h11016: Data = 4'h4; //> 
    18'h11017: Data = 4'h4; //> 
    18'h11018: Data = 4'h4; //> 
    18'h11019: Data = 4'h6; //[ 
    18'h11020: Data = 4'h3; //- 
    18'h11021: Data = 4'h5; //< 
    18'h11022: Data = 4'h5; //< 
    18'h11023: Data = 4'h5; //< 
    18'h11024: Data = 4'h5; //< 
    18'h11025: Data = 4'h2; //+ 
    18'h11026: Data = 4'h4; //> 
    18'h11027: Data = 4'h6; //[ 
    18'h11028: Data = 4'h5; //< 
    18'h11029: Data = 4'h3; //- 
    18'h11030: Data = 4'h4; //> 
    18'h11031: Data = 4'h3; //- 
    18'h11032: Data = 4'h5; //< 
    18'h11033: Data = 4'h5; //< 
    18'h11034: Data = 4'h5; //< 
    18'h11035: Data = 4'h5; //< 
    18'h11036: Data = 4'h5; //< 
    18'h11037: Data = 4'h5; //< 
    18'h11038: Data = 4'h2; //+ 
    18'h11039: Data = 4'h4; //> 
    18'h11040: Data = 4'h4; //> 
    18'h11041: Data = 4'h4; //> 
    18'h11042: Data = 4'h4; //> 
    18'h11043: Data = 4'h4; //> 
    18'h11044: Data = 4'h4; //> 
    18'h11045: Data = 4'h7; //] 
    18'h11046: Data = 4'h5; //< 
    18'h11047: Data = 4'h6; //[ 
    18'h11048: Data = 4'h3; //- 
    18'h11049: Data = 4'h4; //> 
    18'h11050: Data = 4'h2; //+ 
    18'h11051: Data = 4'h5; //< 
    18'h11052: Data = 4'h7; //] 
    18'h11053: Data = 4'h4; //> 
    18'h11054: Data = 4'h4; //> 
    18'h11055: Data = 4'h4; //> 
    18'h11056: Data = 4'h4; //> 
    18'h11057: Data = 4'h7; //] 
    18'h11058: Data = 4'h5; //< 
    18'h11059: Data = 4'h5; //< 
    18'h11060: Data = 4'h5; //< 
    18'h11061: Data = 4'h6; //[ 
    18'h11062: Data = 4'h3; //- 
    18'h11063: Data = 4'h4; //> 
    18'h11064: Data = 4'h4; //> 
    18'h11065: Data = 4'h4; //> 
    18'h11066: Data = 4'h2; //+ 
    18'h11067: Data = 4'h5; //< 
    18'h11068: Data = 4'h5; //< 
    18'h11069: Data = 4'h5; //< 
    18'h11070: Data = 4'h7; //] 
    18'h11071: Data = 4'h5; //< 
    18'h11072: Data = 4'h2; //+ 
    18'h11073: Data = 4'h5; //< 
    18'h11074: Data = 4'h5; //< 
    18'h11075: Data = 4'h5; //< 
    18'h11076: Data = 4'h5; //< 
    18'h11077: Data = 4'h5; //< 
    18'h11078: Data = 4'h5; //< 
    18'h11079: Data = 4'h5; //< 
    18'h11080: Data = 4'h5; //< 
    18'h11081: Data = 4'h5; //< 
    18'h11082: Data = 4'h7; //] 
    18'h11083: Data = 4'h4; //> 
    18'h11084: Data = 4'h4; //> 
    18'h11085: Data = 4'h4; //> 
    18'h11086: Data = 4'h4; //> 
    18'h11087: Data = 4'h4; //> 
    18'h11088: Data = 4'h4; //> 
    18'h11089: Data = 4'h4; //> 
    18'h11090: Data = 4'h4; //> 
    18'h11091: Data = 4'h4; //> 
    18'h11092: Data = 4'h6; //[ 
    18'h11093: Data = 4'h4; //> 
    18'h11094: Data = 4'h2; //+ 
    18'h11095: Data = 4'h4; //> 
    18'h11096: Data = 4'h4; //> 
    18'h11097: Data = 4'h4; //> 
    18'h11098: Data = 4'h4; //> 
    18'h11099: Data = 4'h4; //> 
    18'h11100: Data = 4'h4; //> 
    18'h11101: Data = 4'h4; //> 
    18'h11102: Data = 4'h4; //> 
    18'h11103: Data = 4'h7; //] 
    18'h11104: Data = 4'h5; //< 
    18'h11105: Data = 4'h5; //< 
    18'h11106: Data = 4'h5; //< 
    18'h11107: Data = 4'h5; //< 
    18'h11108: Data = 4'h5; //< 
    18'h11109: Data = 4'h5; //< 
    18'h11110: Data = 4'h5; //< 
    18'h11111: Data = 4'h5; //< 
    18'h11112: Data = 4'h5; //< 
    18'h11113: Data = 4'h6; //[ 
    18'h11114: Data = 4'h5; //< 
    18'h11115: Data = 4'h5; //< 
    18'h11116: Data = 4'h5; //< 
    18'h11117: Data = 4'h5; //< 
    18'h11118: Data = 4'h5; //< 
    18'h11119: Data = 4'h5; //< 
    18'h11120: Data = 4'h5; //< 
    18'h11121: Data = 4'h5; //< 
    18'h11122: Data = 4'h5; //< 
    18'h11123: Data = 4'h7; //] 
    18'h11124: Data = 4'h4; //> 
    18'h11125: Data = 4'h4; //> 
    18'h11126: Data = 4'h4; //> 
    18'h11127: Data = 4'h4; //> 
    18'h11128: Data = 4'h4; //> 
    18'h11129: Data = 4'h4; //> 
    18'h11130: Data = 4'h4; //> 
    18'h11131: Data = 4'h4; //> 
    18'h11132: Data = 4'h4; //> 
    18'h11133: Data = 4'h6; //[ 
    18'h11134: Data = 4'h4; //> 
    18'h11135: Data = 4'h3; //- 
    18'h11136: Data = 4'h4; //> 
    18'h11137: Data = 4'h4; //> 
    18'h11138: Data = 4'h4; //> 
    18'h11139: Data = 4'h4; //> 
    18'h11140: Data = 4'h4; //> 
    18'h11141: Data = 4'h6; //[ 
    18'h11142: Data = 4'h3; //- 
    18'h11143: Data = 4'h5; //< 
    18'h11144: Data = 4'h5; //< 
    18'h11145: Data = 4'h5; //< 
    18'h11146: Data = 4'h5; //< 
    18'h11147: Data = 4'h5; //< 
    18'h11148: Data = 4'h2; //+ 
    18'h11149: Data = 4'h4; //> 
    18'h11150: Data = 4'h4; //> 
    18'h11151: Data = 4'h4; //> 
    18'h11152: Data = 4'h4; //> 
    18'h11153: Data = 4'h4; //> 
    18'h11154: Data = 4'h7; //] 
    18'h11155: Data = 4'h5; //< 
    18'h11156: Data = 4'h5; //< 
    18'h11157: Data = 4'h5; //< 
    18'h11158: Data = 4'h5; //< 
    18'h11159: Data = 4'h5; //< 
    18'h11160: Data = 4'h6; //[ 
    18'h11161: Data = 4'h3; //- 
    18'h11162: Data = 4'h4; //> 
    18'h11163: Data = 4'h4; //> 
    18'h11164: Data = 4'h4; //> 
    18'h11165: Data = 4'h4; //> 
    18'h11166: Data = 4'h4; //> 
    18'h11167: Data = 4'h2; //+ 
    18'h11168: Data = 4'h5; //< 
    18'h11169: Data = 4'h5; //< 
    18'h11170: Data = 4'h5; //< 
    18'h11171: Data = 4'h5; //< 
    18'h11172: Data = 4'h5; //< 
    18'h11173: Data = 4'h5; //< 
    18'h11174: Data = 4'h6; //[ 
    18'h11175: Data = 4'h3; //- 
    18'h11176: Data = 4'h4; //> 
    18'h11177: Data = 4'h4; //> 
    18'h11178: Data = 4'h4; //> 
    18'h11179: Data = 4'h6; //[ 
    18'h11180: Data = 4'h3; //- 
    18'h11181: Data = 4'h5; //< 
    18'h11182: Data = 4'h5; //< 
    18'h11183: Data = 4'h5; //< 
    18'h11184: Data = 4'h2; //+ 
    18'h11185: Data = 4'h4; //> 
    18'h11186: Data = 4'h4; //> 
    18'h11187: Data = 4'h4; //> 
    18'h11188: Data = 4'h7; //] 
    18'h11189: Data = 4'h5; //< 
    18'h11190: Data = 4'h5; //< 
    18'h11191: Data = 4'h5; //< 
    18'h11192: Data = 4'h6; //[ 
    18'h11193: Data = 4'h3; //- 
    18'h11194: Data = 4'h4; //> 
    18'h11195: Data = 4'h4; //> 
    18'h11196: Data = 4'h4; //> 
    18'h11197: Data = 4'h2; //+ 
    18'h11198: Data = 4'h4; //> 
    18'h11199: Data = 4'h2; //+ 
    18'h11200: Data = 4'h5; //< 
    18'h11201: Data = 4'h5; //< 
    18'h11202: Data = 4'h5; //< 
    18'h11203: Data = 4'h5; //< 
    18'h11204: Data = 4'h7; //] 
    18'h11205: Data = 4'h2; //+ 
    18'h11206: Data = 4'h4; //> 
    18'h11207: Data = 4'h4; //> 
    18'h11208: Data = 4'h4; //> 
    18'h11209: Data = 4'h4; //> 
    18'h11210: Data = 4'h4; //> 
    18'h11211: Data = 4'h4; //> 
    18'h11212: Data = 4'h4; //> 
    18'h11213: Data = 4'h4; //> 
    18'h11214: Data = 4'h4; //> 
    18'h11215: Data = 4'h7; //] 
    18'h11216: Data = 4'h5; //< 
    18'h11217: Data = 4'h5; //< 
    18'h11218: Data = 4'h5; //< 
    18'h11219: Data = 4'h5; //< 
    18'h11220: Data = 4'h5; //< 
    18'h11221: Data = 4'h5; //< 
    18'h11222: Data = 4'h5; //< 
    18'h11223: Data = 4'h5; //< 
    18'h11224: Data = 4'h6; //[ 
    18'h11225: Data = 4'h5; //< 
    18'h11226: Data = 4'h5; //< 
    18'h11227: Data = 4'h5; //< 
    18'h11228: Data = 4'h5; //< 
    18'h11229: Data = 4'h5; //< 
    18'h11230: Data = 4'h5; //< 
    18'h11231: Data = 4'h5; //< 
    18'h11232: Data = 4'h5; //< 
    18'h11233: Data = 4'h5; //< 
    18'h11234: Data = 4'h7; //] 
    18'h11235: Data = 4'h7; //] 
    18'h11236: Data = 4'h4; //> 
    18'h11237: Data = 4'h4; //> 
    18'h11238: Data = 4'h4; //> 
    18'h11239: Data = 4'h4; //> 
    18'h11240: Data = 4'h4; //> 
    18'h11241: Data = 4'h4; //> 
    18'h11242: Data = 4'h4; //> 
    18'h11243: Data = 4'h4; //> 
    18'h11244: Data = 4'h4; //> 
    18'h11245: Data = 4'h6; //[ 
    18'h11246: Data = 4'h4; //> 
    18'h11247: Data = 4'h4; //> 
    18'h11248: Data = 4'h4; //> 
    18'h11249: Data = 4'h4; //> 
    18'h11250: Data = 4'h4; //> 
    18'h11251: Data = 4'h4; //> 
    18'h11252: Data = 4'h4; //> 
    18'h11253: Data = 4'h4; //> 
    18'h11254: Data = 4'h4; //> 
    18'h11255: Data = 4'h7; //] 
    18'h11256: Data = 4'h5; //< 
    18'h11257: Data = 4'h5; //< 
    18'h11258: Data = 4'h5; //< 
    18'h11259: Data = 4'h5; //< 
    18'h11260: Data = 4'h5; //< 
    18'h11261: Data = 4'h5; //< 
    18'h11262: Data = 4'h5; //< 
    18'h11263: Data = 4'h5; //< 
    18'h11264: Data = 4'h5; //< 
    18'h11265: Data = 4'h6; //[ 
    18'h11266: Data = 4'h4; //> 
    18'h11267: Data = 4'h4; //> 
    18'h11268: Data = 4'h6; //[ 
    18'h11269: Data = 4'h3; //- 
    18'h11270: Data = 4'h4; //> 
    18'h11271: Data = 4'h4; //> 
    18'h11272: Data = 4'h4; //> 
    18'h11273: Data = 4'h4; //> 
    18'h11274: Data = 4'h4; //> 
    18'h11275: Data = 4'h4; //> 
    18'h11276: Data = 4'h4; //> 
    18'h11277: Data = 4'h4; //> 
    18'h11278: Data = 4'h4; //> 
    18'h11279: Data = 4'h2; //+ 
    18'h11280: Data = 4'h5; //< 
    18'h11281: Data = 4'h5; //< 
    18'h11282: Data = 4'h5; //< 
    18'h11283: Data = 4'h5; //< 
    18'h11284: Data = 4'h5; //< 
    18'h11285: Data = 4'h5; //< 
    18'h11286: Data = 4'h5; //< 
    18'h11287: Data = 4'h5; //< 
    18'h11288: Data = 4'h5; //< 
    18'h11289: Data = 4'h7; //] 
    18'h11290: Data = 4'h5; //< 
    18'h11291: Data = 4'h5; //< 
    18'h11292: Data = 4'h5; //< 
    18'h11293: Data = 4'h5; //< 
    18'h11294: Data = 4'h5; //< 
    18'h11295: Data = 4'h5; //< 
    18'h11296: Data = 4'h5; //< 
    18'h11297: Data = 4'h5; //< 
    18'h11298: Data = 4'h5; //< 
    18'h11299: Data = 4'h5; //< 
    18'h11300: Data = 4'h5; //< 
    18'h11301: Data = 4'h7; //] 
    18'h11302: Data = 4'h4; //> 
    18'h11303: Data = 4'h4; //> 
    18'h11304: Data = 4'h6; //[ 
    18'h11305: Data = 4'h3; //- 
    18'h11306: Data = 4'h4; //> 
    18'h11307: Data = 4'h4; //> 
    18'h11308: Data = 4'h4; //> 
    18'h11309: Data = 4'h4; //> 
    18'h11310: Data = 4'h4; //> 
    18'h11311: Data = 4'h4; //> 
    18'h11312: Data = 4'h4; //> 
    18'h11313: Data = 4'h4; //> 
    18'h11314: Data = 4'h4; //> 
    18'h11315: Data = 4'h2; //+ 
    18'h11316: Data = 4'h5; //< 
    18'h11317: Data = 4'h5; //< 
    18'h11318: Data = 4'h5; //< 
    18'h11319: Data = 4'h5; //< 
    18'h11320: Data = 4'h5; //< 
    18'h11321: Data = 4'h5; //< 
    18'h11322: Data = 4'h5; //< 
    18'h11323: Data = 4'h5; //< 
    18'h11324: Data = 4'h5; //< 
    18'h11325: Data = 4'h7; //] 
    18'h11326: Data = 4'h5; //< 
    18'h11327: Data = 4'h5; //< 
    18'h11328: Data = 4'h2; //+ 
    18'h11329: Data = 4'h4; //> 
    18'h11330: Data = 4'h4; //> 
    18'h11331: Data = 4'h4; //> 
    18'h11332: Data = 4'h4; //> 
    18'h11333: Data = 4'h4; //> 
    18'h11334: Data = 4'h4; //> 
    18'h11335: Data = 4'h4; //> 
    18'h11336: Data = 4'h4; //> 
    18'h11337: Data = 4'h7; //] 
    18'h11338: Data = 4'h5; //< 
    18'h11339: Data = 4'h5; //< 
    18'h11340: Data = 4'h5; //< 
    18'h11341: Data = 4'h5; //< 
    18'h11342: Data = 4'h5; //< 
    18'h11343: Data = 4'h5; //< 
    18'h11344: Data = 4'h5; //< 
    18'h11345: Data = 4'h5; //< 
    18'h11346: Data = 4'h5; //< 
    18'h11347: Data = 4'h6; //[ 
    18'h11348: Data = 4'h4; //> 
    18'h11349: Data = 4'ha; //0 
    18'h11350: Data = 4'h5; //< 
    18'h11351: Data = 4'h3; //- 
    18'h11352: Data = 4'h4; //> 
    18'h11353: Data = 4'h4; //> 
    18'h11354: Data = 4'h4; //> 
    18'h11355: Data = 4'h4; //> 
    18'h11356: Data = 4'h6; //[ 
    18'h11357: Data = 4'h3; //- 
    18'h11358: Data = 4'h5; //< 
    18'h11359: Data = 4'h5; //< 
    18'h11360: Data = 4'h5; //< 
    18'h11361: Data = 4'h5; //< 
    18'h11362: Data = 4'h2; //+ 
    18'h11363: Data = 4'h4; //> 
    18'h11364: Data = 4'h6; //[ 
    18'h11365: Data = 4'h5; //< 
    18'h11366: Data = 4'h3; //- 
    18'h11367: Data = 4'h4; //> 
    18'h11368: Data = 4'h3; //- 
    18'h11369: Data = 4'h5; //< 
    18'h11370: Data = 4'h5; //< 
    18'h11371: Data = 4'h5; //< 
    18'h11372: Data = 4'h5; //< 
    18'h11373: Data = 4'h5; //< 
    18'h11374: Data = 4'h5; //< 
    18'h11375: Data = 4'h2; //+ 
    18'h11376: Data = 4'h4; //> 
    18'h11377: Data = 4'h4; //> 
    18'h11378: Data = 4'h4; //> 
    18'h11379: Data = 4'h4; //> 
    18'h11380: Data = 4'h4; //> 
    18'h11381: Data = 4'h4; //> 
    18'h11382: Data = 4'h7; //] 
    18'h11383: Data = 4'h5; //< 
    18'h11384: Data = 4'h6; //[ 
    18'h11385: Data = 4'h3; //- 
    18'h11386: Data = 4'h4; //> 
    18'h11387: Data = 4'h2; //+ 
    18'h11388: Data = 4'h5; //< 
    18'h11389: Data = 4'h7; //] 
    18'h11390: Data = 4'h4; //> 
    18'h11391: Data = 4'h4; //> 
    18'h11392: Data = 4'h4; //> 
    18'h11393: Data = 4'h4; //> 
    18'h11394: Data = 4'h7; //] 
    18'h11395: Data = 4'h5; //< 
    18'h11396: Data = 4'h5; //< 
    18'h11397: Data = 4'h5; //< 
    18'h11398: Data = 4'h6; //[ 
    18'h11399: Data = 4'h3; //- 
    18'h11400: Data = 4'h4; //> 
    18'h11401: Data = 4'h4; //> 
    18'h11402: Data = 4'h4; //> 
    18'h11403: Data = 4'h2; //+ 
    18'h11404: Data = 4'h5; //< 
    18'h11405: Data = 4'h5; //< 
    18'h11406: Data = 4'h5; //< 
    18'h11407: Data = 4'h7; //] 
    18'h11408: Data = 4'h5; //< 
    18'h11409: Data = 4'h2; //+ 
    18'h11410: Data = 4'h5; //< 
    18'h11411: Data = 4'h5; //< 
    18'h11412: Data = 4'h5; //< 
    18'h11413: Data = 4'h5; //< 
    18'h11414: Data = 4'h5; //< 
    18'h11415: Data = 4'h5; //< 
    18'h11416: Data = 4'h5; //< 
    18'h11417: Data = 4'h5; //< 
    18'h11418: Data = 4'h5; //< 
    18'h11419: Data = 4'h7; //] 
    18'h11420: Data = 4'h4; //> 
    18'h11421: Data = 4'h4; //> 
    18'h11422: Data = 4'h4; //> 
    18'h11423: Data = 4'h4; //> 
    18'h11424: Data = 4'h4; //> 
    18'h11425: Data = 4'h4; //> 
    18'h11426: Data = 4'h4; //> 
    18'h11427: Data = 4'h4; //> 
    18'h11428: Data = 4'h4; //> 
    18'h11429: Data = 4'h6; //[ 
    18'h11430: Data = 4'h4; //> 
    18'h11431: Data = 4'h4; //> 
    18'h11432: Data = 4'h4; //> 
    18'h11433: Data = 4'h4; //> 
    18'h11434: Data = 4'h6; //[ 
    18'h11435: Data = 4'h3; //- 
    18'h11436: Data = 4'h5; //< 
    18'h11437: Data = 4'h5; //< 
    18'h11438: Data = 4'h5; //< 
    18'h11439: Data = 4'h5; //< 
    18'h11440: Data = 4'h5; //< 
    18'h11441: Data = 4'h5; //< 
    18'h11442: Data = 4'h5; //< 
    18'h11443: Data = 4'h5; //< 
    18'h11444: Data = 4'h5; //< 
    18'h11445: Data = 4'h5; //< 
    18'h11446: Data = 4'h5; //< 
    18'h11447: Data = 4'h5; //< 
    18'h11448: Data = 4'h5; //< 
    18'h11449: Data = 4'h5; //< 
    18'h11450: Data = 4'h5; //< 
    18'h11451: Data = 4'h5; //< 
    18'h11452: Data = 4'h5; //< 
    18'h11453: Data = 4'h5; //< 
    18'h11454: Data = 4'h5; //< 
    18'h11455: Data = 4'h5; //< 
    18'h11456: Data = 4'h5; //< 
    18'h11457: Data = 4'h5; //< 
    18'h11458: Data = 4'h5; //< 
    18'h11459: Data = 4'h5; //< 
    18'h11460: Data = 4'h5; //< 
    18'h11461: Data = 4'h5; //< 
    18'h11462: Data = 4'h5; //< 
    18'h11463: Data = 4'h5; //< 
    18'h11464: Data = 4'h5; //< 
    18'h11465: Data = 4'h5; //< 
    18'h11466: Data = 4'h5; //< 
    18'h11467: Data = 4'h5; //< 
    18'h11468: Data = 4'h5; //< 
    18'h11469: Data = 4'h5; //< 
    18'h11470: Data = 4'h5; //< 
    18'h11471: Data = 4'h5; //< 
    18'h11472: Data = 4'h2; //+ 
    18'h11473: Data = 4'h4; //> 
    18'h11474: Data = 4'h4; //> 
    18'h11475: Data = 4'h4; //> 
    18'h11476: Data = 4'h4; //> 
    18'h11477: Data = 4'h4; //> 
    18'h11478: Data = 4'h4; //> 
    18'h11479: Data = 4'h4; //> 
    18'h11480: Data = 4'h4; //> 
    18'h11481: Data = 4'h4; //> 
    18'h11482: Data = 4'h4; //> 
    18'h11483: Data = 4'h4; //> 
    18'h11484: Data = 4'h4; //> 
    18'h11485: Data = 4'h4; //> 
    18'h11486: Data = 4'h4; //> 
    18'h11487: Data = 4'h4; //> 
    18'h11488: Data = 4'h4; //> 
    18'h11489: Data = 4'h4; //> 
    18'h11490: Data = 4'h4; //> 
    18'h11491: Data = 4'h4; //> 
    18'h11492: Data = 4'h4; //> 
    18'h11493: Data = 4'h4; //> 
    18'h11494: Data = 4'h4; //> 
    18'h11495: Data = 4'h4; //> 
    18'h11496: Data = 4'h4; //> 
    18'h11497: Data = 4'h4; //> 
    18'h11498: Data = 4'h4; //> 
    18'h11499: Data = 4'h4; //> 
    18'h11500: Data = 4'h4; //> 
    18'h11501: Data = 4'h4; //> 
    18'h11502: Data = 4'h4; //> 
    18'h11503: Data = 4'h4; //> 
    18'h11504: Data = 4'h4; //> 
    18'h11505: Data = 4'h4; //> 
    18'h11506: Data = 4'h4; //> 
    18'h11507: Data = 4'h4; //> 
    18'h11508: Data = 4'h4; //> 
    18'h11509: Data = 4'h7; //] 
    18'h11510: Data = 4'h4; //> 
    18'h11511: Data = 4'h4; //> 
    18'h11512: Data = 4'h4; //> 
    18'h11513: Data = 4'h4; //> 
    18'h11514: Data = 4'h4; //> 
    18'h11515: Data = 4'h7; //] 
    18'h11516: Data = 4'h5; //< 
    18'h11517: Data = 4'h5; //< 
    18'h11518: Data = 4'h5; //< 
    18'h11519: Data = 4'h5; //< 
    18'h11520: Data = 4'h5; //< 
    18'h11521: Data = 4'h5; //< 
    18'h11522: Data = 4'h5; //< 
    18'h11523: Data = 4'h5; //< 
    18'h11524: Data = 4'h5; //< 
    18'h11525: Data = 4'h6; //[ 
    18'h11526: Data = 4'h5; //< 
    18'h11527: Data = 4'h5; //< 
    18'h11528: Data = 4'h5; //< 
    18'h11529: Data = 4'h5; //< 
    18'h11530: Data = 4'h5; //< 
    18'h11531: Data = 4'h5; //< 
    18'h11532: Data = 4'h5; //< 
    18'h11533: Data = 4'h5; //< 
    18'h11534: Data = 4'h5; //< 
    18'h11535: Data = 4'h7; //] 
    18'h11536: Data = 4'h4; //> 
    18'h11537: Data = 4'h4; //> 
    18'h11538: Data = 4'h4; //> 
    18'h11539: Data = 4'h4; //> 
    18'h11540: Data = 4'h4; //> 
    18'h11541: Data = 4'h4; //> 
    18'h11542: Data = 4'h4; //> 
    18'h11543: Data = 4'h4; //> 
    18'h11544: Data = 4'h4; //> 
    18'h11545: Data = 4'h2; //+ 
    18'h11546: Data = 4'h2; //+ 
    18'h11547: Data = 4'h2; //+ 
    18'h11548: Data = 4'h2; //+ 
    18'h11549: Data = 4'h2; //+ 
    18'h11550: Data = 4'h2; //+ 
    18'h11551: Data = 4'h2; //+ 
    18'h11552: Data = 4'h2; //+ 
    18'h11553: Data = 4'h2; //+ 
    18'h11554: Data = 4'h2; //+ 
    18'h11555: Data = 4'h2; //+ 
    18'h11556: Data = 4'h2; //+ 
    18'h11557: Data = 4'h2; //+ 
    18'h11558: Data = 4'h2; //+ 
    18'h11559: Data = 4'h2; //+ 
    18'h11560: Data = 4'h6; //[ 
    18'h11561: Data = 4'h6; //[ 
    18'h11562: Data = 4'h4; //> 
    18'h11563: Data = 4'h4; //> 
    18'h11564: Data = 4'h4; //> 
    18'h11565: Data = 4'h4; //> 
    18'h11566: Data = 4'h4; //> 
    18'h11567: Data = 4'h4; //> 
    18'h11568: Data = 4'h4; //> 
    18'h11569: Data = 4'h4; //> 
    18'h11570: Data = 4'h4; //> 
    18'h11571: Data = 4'h7; //] 
    18'h11572: Data = 4'h5; //< 
    18'h11573: Data = 4'h5; //< 
    18'h11574: Data = 4'h5; //< 
    18'h11575: Data = 4'h5; //< 
    18'h11576: Data = 4'h5; //< 
    18'h11577: Data = 4'h5; //< 
    18'h11578: Data = 4'h5; //< 
    18'h11579: Data = 4'h5; //< 
    18'h11580: Data = 4'h5; //< 
    18'h11581: Data = 4'h3; //- 
    18'h11582: Data = 4'h5; //< 
    18'h11583: Data = 4'h5; //< 
    18'h11584: Data = 4'h5; //< 
    18'h11585: Data = 4'h5; //< 
    18'h11586: Data = 4'h5; //< 
    18'h11587: Data = 4'h5; //< 
    18'h11588: Data = 4'h5; //< 
    18'h11589: Data = 4'h5; //< 
    18'h11590: Data = 4'h5; //< 
    18'h11591: Data = 4'h6; //[ 
    18'h11592: Data = 4'h5; //< 
    18'h11593: Data = 4'h5; //< 
    18'h11594: Data = 4'h5; //< 
    18'h11595: Data = 4'h5; //< 
    18'h11596: Data = 4'h5; //< 
    18'h11597: Data = 4'h5; //< 
    18'h11598: Data = 4'h5; //< 
    18'h11599: Data = 4'h5; //< 
    18'h11600: Data = 4'h5; //< 
    18'h11601: Data = 4'h7; //] 
    18'h11602: Data = 4'h4; //> 
    18'h11603: Data = 4'h4; //> 
    18'h11604: Data = 4'h4; //> 
    18'h11605: Data = 4'h4; //> 
    18'h11606: Data = 4'h4; //> 
    18'h11607: Data = 4'h4; //> 
    18'h11608: Data = 4'h4; //> 
    18'h11609: Data = 4'h4; //> 
    18'h11610: Data = 4'h4; //> 
    18'h11611: Data = 4'h3; //- 
    18'h11612: Data = 4'h7; //] 
    18'h11613: Data = 4'h2; //+ 
    18'h11614: Data = 4'h4; //> 
    18'h11615: Data = 4'h4; //> 
    18'h11616: Data = 4'h4; //> 
    18'h11617: Data = 4'h4; //> 
    18'h11618: Data = 4'h4; //> 
    18'h11619: Data = 4'h4; //> 
    18'h11620: Data = 4'h4; //> 
    18'h11621: Data = 4'h4; //> 
    18'h11622: Data = 4'h4; //> 
    18'h11623: Data = 4'h4; //> 
    18'h11624: Data = 4'h4; //> 
    18'h11625: Data = 4'h4; //> 
    18'h11626: Data = 4'h4; //> 
    18'h11627: Data = 4'h4; //> 
    18'h11628: Data = 4'h4; //> 
    18'h11629: Data = 4'h4; //> 
    18'h11630: Data = 4'h4; //> 
    18'h11631: Data = 4'h4; //> 
    18'h11632: Data = 4'h4; //> 
    18'h11633: Data = 4'h4; //> 
    18'h11634: Data = 4'h4; //> 
    18'h11635: Data = 4'h2; //+ 
    18'h11636: Data = 4'h5; //< 
    18'h11637: Data = 4'h5; //< 
    18'h11638: Data = 4'h5; //< 
    18'h11639: Data = 4'h6; //[ 
    18'h11640: Data = 4'h5; //< 
    18'h11641: Data = 4'h5; //< 
    18'h11642: Data = 4'h5; //< 
    18'h11643: Data = 4'h5; //< 
    18'h11644: Data = 4'h5; //< 
    18'h11645: Data = 4'h5; //< 
    18'h11646: Data = 4'h5; //< 
    18'h11647: Data = 4'h5; //< 
    18'h11648: Data = 4'h5; //< 
    18'h11649: Data = 4'h7; //] 
    18'h11650: Data = 4'h4; //> 
    18'h11651: Data = 4'h4; //> 
    18'h11652: Data = 4'h4; //> 
    18'h11653: Data = 4'h4; //> 
    18'h11654: Data = 4'h4; //> 
    18'h11655: Data = 4'h4; //> 
    18'h11656: Data = 4'h4; //> 
    18'h11657: Data = 4'h4; //> 
    18'h11658: Data = 4'h4; //> 
    18'h11659: Data = 4'h6; //[ 
    18'h11660: Data = 4'h4; //> 
    18'h11661: Data = 4'h4; //> 
    18'h11662: Data = 4'h4; //> 
    18'h11663: Data = 4'h6; //[ 
    18'h11664: Data = 4'h3; //- 
    18'h11665: Data = 4'h5; //< 
    18'h11666: Data = 4'h5; //< 
    18'h11667: Data = 4'h5; //< 
    18'h11668: Data = 4'h3; //- 
    18'h11669: Data = 4'h4; //> 
    18'h11670: Data = 4'h4; //> 
    18'h11671: Data = 4'h4; //> 
    18'h11672: Data = 4'h7; //] 
    18'h11673: Data = 4'h2; //+ 
    18'h11674: Data = 4'h5; //< 
    18'h11675: Data = 4'h5; //< 
    18'h11676: Data = 4'h5; //< 
    18'h11677: Data = 4'h6; //[ 
    18'h11678: Data = 4'h3; //- 
    18'h11679: Data = 4'h4; //> 
    18'h11680: Data = 4'h4; //> 
    18'h11681: Data = 4'h4; //> 
    18'h11682: Data = 4'h3; //- 
    18'h11683: Data = 4'h4; //> 
    18'h11684: Data = 4'h6; //[ 
    18'h11685: Data = 4'h3; //- 
    18'h11686: Data = 4'h5; //< 
    18'h11687: Data = 4'h5; //< 
    18'h11688: Data = 4'h5; //< 
    18'h11689: Data = 4'h5; //< 
    18'h11690: Data = 4'h2; //+ 
    18'h11691: Data = 4'h4; //> 
    18'h11692: Data = 4'h4; //> 
    18'h11693: Data = 4'h4; //> 
    18'h11694: Data = 4'h4; //> 
    18'h11695: Data = 4'h7; //] 
    18'h11696: Data = 4'h5; //< 
    18'h11697: Data = 4'h5; //< 
    18'h11698: Data = 4'h5; //< 
    18'h11699: Data = 4'h5; //< 
    18'h11700: Data = 4'h6; //[ 
    18'h11701: Data = 4'h3; //- 
    18'h11702: Data = 4'h4; //> 
    18'h11703: Data = 4'h4; //> 
    18'h11704: Data = 4'h4; //> 
    18'h11705: Data = 4'h4; //> 
    18'h11706: Data = 4'h2; //+ 
    18'h11707: Data = 4'h5; //< 
    18'h11708: Data = 4'h5; //< 
    18'h11709: Data = 4'h5; //< 
    18'h11710: Data = 4'h5; //< 
    18'h11711: Data = 4'h5; //< 
    18'h11712: Data = 4'h5; //< 
    18'h11713: Data = 4'h5; //< 
    18'h11714: Data = 4'h5; //< 
    18'h11715: Data = 4'h5; //< 
    18'h11716: Data = 4'h5; //< 
    18'h11717: Data = 4'h5; //< 
    18'h11718: Data = 4'h5; //< 
    18'h11719: Data = 4'h5; //< 
    18'h11720: Data = 4'h6; //[ 
    18'h11721: Data = 4'h5; //< 
    18'h11722: Data = 4'h5; //< 
    18'h11723: Data = 4'h5; //< 
    18'h11724: Data = 4'h5; //< 
    18'h11725: Data = 4'h5; //< 
    18'h11726: Data = 4'h5; //< 
    18'h11727: Data = 4'h5; //< 
    18'h11728: Data = 4'h5; //< 
    18'h11729: Data = 4'h5; //< 
    18'h11730: Data = 4'h7; //] 
    18'h11731: Data = 4'h4; //> 
    18'h11732: Data = 4'h4; //> 
    18'h11733: Data = 4'h4; //> 
    18'h11734: Data = 4'h4; //> 
    18'h11735: Data = 4'ha; //0 
    18'h11736: Data = 4'h2; //+ 
    18'h11737: Data = 4'h4; //> 
    18'h11738: Data = 4'h4; //> 
    18'h11739: Data = 4'h4; //> 
    18'h11740: Data = 4'h4; //> 
    18'h11741: Data = 4'h4; //> 
    18'h11742: Data = 4'h6; //[ 
    18'h11743: Data = 4'h4; //> 
    18'h11744: Data = 4'h4; //> 
    18'h11745: Data = 4'h4; //> 
    18'h11746: Data = 4'h4; //> 
    18'h11747: Data = 4'h4; //> 
    18'h11748: Data = 4'h4; //> 
    18'h11749: Data = 4'h4; //> 
    18'h11750: Data = 4'h4; //> 
    18'h11751: Data = 4'h4; //> 
    18'h11752: Data = 4'h7; //] 
    18'h11753: Data = 4'h4; //> 
    18'h11754: Data = 4'h2; //+ 
    18'h11755: Data = 4'h5; //< 
    18'h11756: Data = 4'h7; //] 
    18'h11757: Data = 4'h7; //] 
    18'h11758: Data = 4'h2; //+ 
    18'h11759: Data = 4'h4; //> 
    18'h11760: Data = 4'h4; //> 
    18'h11761: Data = 4'h4; //> 
    18'h11762: Data = 4'h4; //> 
    18'h11763: Data = 4'h6; //[ 
    18'h11764: Data = 4'h3; //- 
    18'h11765: Data = 4'h5; //< 
    18'h11766: Data = 4'h5; //< 
    18'h11767: Data = 4'h5; //< 
    18'h11768: Data = 4'h5; //< 
    18'h11769: Data = 4'h3; //- 
    18'h11770: Data = 4'h4; //> 
    18'h11771: Data = 4'h4; //> 
    18'h11772: Data = 4'h4; //> 
    18'h11773: Data = 4'h4; //> 
    18'h11774: Data = 4'h7; //] 
    18'h11775: Data = 4'h2; //+ 
    18'h11776: Data = 4'h5; //< 
    18'h11777: Data = 4'h5; //< 
    18'h11778: Data = 4'h5; //< 
    18'h11779: Data = 4'h5; //< 
    18'h11780: Data = 4'h6; //[ 
    18'h11781: Data = 4'h3; //- 
    18'h11782: Data = 4'h4; //> 
    18'h11783: Data = 4'h4; //> 
    18'h11784: Data = 4'h4; //> 
    18'h11785: Data = 4'h4; //> 
    18'h11786: Data = 4'h3; //- 
    18'h11787: Data = 4'h5; //< 
    18'h11788: Data = 4'h6; //[ 
    18'h11789: Data = 4'h3; //- 
    18'h11790: Data = 4'h5; //< 
    18'h11791: Data = 4'h5; //< 
    18'h11792: Data = 4'h5; //< 
    18'h11793: Data = 4'h2; //+ 
    18'h11794: Data = 4'h4; //> 
    18'h11795: Data = 4'h4; //> 
    18'h11796: Data = 4'h4; //> 
    18'h11797: Data = 4'h7; //] 
    18'h11798: Data = 4'h5; //< 
    18'h11799: Data = 4'h5; //< 
    18'h11800: Data = 4'h5; //< 
    18'h11801: Data = 4'h6; //[ 
    18'h11802: Data = 4'h3; //- 
    18'h11803: Data = 4'h4; //> 
    18'h11804: Data = 4'h4; //> 
    18'h11805: Data = 4'h4; //> 
    18'h11806: Data = 4'h2; //+ 
    18'h11807: Data = 4'h5; //< 
    18'h11808: Data = 4'h5; //< 
    18'h11809: Data = 4'h5; //< 
    18'h11810: Data = 4'h5; //< 
    18'h11811: Data = 4'h5; //< 
    18'h11812: Data = 4'h5; //< 
    18'h11813: Data = 4'h5; //< 
    18'h11814: Data = 4'h5; //< 
    18'h11815: Data = 4'h5; //< 
    18'h11816: Data = 4'h5; //< 
    18'h11817: Data = 4'h5; //< 
    18'h11818: Data = 4'h5; //< 
    18'h11819: Data = 4'h6; //[ 
    18'h11820: Data = 4'h5; //< 
    18'h11821: Data = 4'h5; //< 
    18'h11822: Data = 4'h5; //< 
    18'h11823: Data = 4'h5; //< 
    18'h11824: Data = 4'h5; //< 
    18'h11825: Data = 4'h5; //< 
    18'h11826: Data = 4'h5; //< 
    18'h11827: Data = 4'h5; //< 
    18'h11828: Data = 4'h5; //< 
    18'h11829: Data = 4'h7; //] 
    18'h11830: Data = 4'h4; //> 
    18'h11831: Data = 4'h4; //> 
    18'h11832: Data = 4'h4; //> 
    18'h11833: Data = 4'ha; //0 
    18'h11834: Data = 4'h2; //+ 
    18'h11835: Data = 4'h4; //> 
    18'h11836: Data = 4'h4; //> 
    18'h11837: Data = 4'h4; //> 
    18'h11838: Data = 4'h4; //> 
    18'h11839: Data = 4'h4; //> 
    18'h11840: Data = 4'h4; //> 
    18'h11841: Data = 4'h6; //[ 
    18'h11842: Data = 4'h4; //> 
    18'h11843: Data = 4'h4; //> 
    18'h11844: Data = 4'h4; //> 
    18'h11845: Data = 4'h4; //> 
    18'h11846: Data = 4'h4; //> 
    18'h11847: Data = 4'h4; //> 
    18'h11848: Data = 4'h4; //> 
    18'h11849: Data = 4'h4; //> 
    18'h11850: Data = 4'h4; //> 
    18'h11851: Data = 4'h7; //] 
    18'h11852: Data = 4'h4; //> 
    18'h11853: Data = 4'ha; //0 
    18'h11854: Data = 4'h2; //+ 
    18'h11855: Data = 4'h5; //< 
    18'h11856: Data = 4'h7; //] 
    18'h11857: Data = 4'h7; //] 
    18'h11858: Data = 4'h2; //+ 
    18'h11859: Data = 4'h4; //> 
    18'h11860: Data = 4'h6; //[ 
    18'h11861: Data = 4'h3; //- 
    18'h11862: Data = 4'h5; //< 
    18'h11863: Data = 4'h6; //[ 
    18'h11864: Data = 4'h4; //> 
    18'h11865: Data = 4'h4; //> 
    18'h11866: Data = 4'h4; //> 
    18'h11867: Data = 4'h4; //> 
    18'h11868: Data = 4'h4; //> 
    18'h11869: Data = 4'h4; //> 
    18'h11870: Data = 4'h4; //> 
    18'h11871: Data = 4'h4; //> 
    18'h11872: Data = 4'h4; //> 
    18'h11873: Data = 4'h7; //] 
    18'h11874: Data = 4'h5; //< 
    18'h11875: Data = 4'h5; //< 
    18'h11876: Data = 4'h5; //< 
    18'h11877: Data = 4'h5; //< 
    18'h11878: Data = 4'h5; //< 
    18'h11879: Data = 4'h5; //< 
    18'h11880: Data = 4'h5; //< 
    18'h11881: Data = 4'h5; //< 
    18'h11882: Data = 4'h7; //] 
    18'h11883: Data = 4'h4; //> 
    18'h11884: Data = 4'h4; //> 
    18'h11885: Data = 4'h4; //> 
    18'h11886: Data = 4'h4; //> 
    18'h11887: Data = 4'h4; //> 
    18'h11888: Data = 4'h4; //> 
    18'h11889: Data = 4'h4; //> 
    18'h11890: Data = 4'h4; //> 
    18'h11891: Data = 4'h7; //] 
    18'h11892: Data = 4'h5; //< 
    18'h11893: Data = 4'h5; //< 
    18'h11894: Data = 4'h5; //< 
    18'h11895: Data = 4'h5; //< 
    18'h11896: Data = 4'h5; //< 
    18'h11897: Data = 4'h5; //< 
    18'h11898: Data = 4'h5; //< 
    18'h11899: Data = 4'h5; //< 
    18'h11900: Data = 4'h5; //< 
    18'h11901: Data = 4'h6; //[ 
    18'h11902: Data = 4'h5; //< 
    18'h11903: Data = 4'h5; //< 
    18'h11904: Data = 4'h5; //< 
    18'h11905: Data = 4'h5; //< 
    18'h11906: Data = 4'h5; //< 
    18'h11907: Data = 4'h5; //< 
    18'h11908: Data = 4'h5; //< 
    18'h11909: Data = 4'h5; //< 
    18'h11910: Data = 4'h5; //< 
    18'h11911: Data = 4'h7; //] 
    18'h11912: Data = 4'h5; //< 
    18'h11913: Data = 4'h5; //< 
    18'h11914: Data = 4'h5; //< 
    18'h11915: Data = 4'h5; //< 
    18'h11916: Data = 4'h5; //< 
    18'h11917: Data = 4'h5; //< 
    18'h11918: Data = 4'h5; //< 
    18'h11919: Data = 4'h6; //[ 
    18'h11920: Data = 4'h3; //- 
    18'h11921: Data = 4'h4; //> 
    18'h11922: Data = 4'h2; //+ 
    18'h11923: Data = 4'h4; //> 
    18'h11924: Data = 4'h4; //> 
    18'h11925: Data = 4'h4; //> 
    18'h11926: Data = 4'h3; //- 
    18'h11927: Data = 4'h5; //< 
    18'h11928: Data = 4'h5; //< 
    18'h11929: Data = 4'h5; //< 
    18'h11930: Data = 4'h5; //< 
    18'h11931: Data = 4'h7; //] 
    18'h11932: Data = 4'h4; //> 
    18'h11933: Data = 4'h4; //> 
    18'h11934: Data = 4'h4; //> 
    18'h11935: Data = 4'h4; //> 
    18'h11936: Data = 4'h4; //> 
    18'h11937: Data = 4'h4; //> 
    18'h11938: Data = 4'h4; //> 
    18'h11939: Data = 4'h4; //> 
    18'h11940: Data = 4'h4; //> 
    18'h11941: Data = 4'h2; //+ 
    18'h11942: Data = 4'h2; //+ 
    18'h11943: Data = 4'h2; //+ 
    18'h11944: Data = 4'h2; //+ 
    18'h11945: Data = 4'h2; //+ 
    18'h11946: Data = 4'h2; //+ 
    18'h11947: Data = 4'h2; //+ 
    18'h11948: Data = 4'h2; //+ 
    18'h11949: Data = 4'h2; //+ 
    18'h11950: Data = 4'h2; //+ 
    18'h11951: Data = 4'h2; //+ 
    18'h11952: Data = 4'h2; //+ 
    18'h11953: Data = 4'h2; //+ 
    18'h11954: Data = 4'h2; //+ 
    18'h11955: Data = 4'h2; //+ 
    18'h11956: Data = 4'h2; //+ 
    18'h11957: Data = 4'h2; //+ 
    18'h11958: Data = 4'h2; //+ 
    18'h11959: Data = 4'h2; //+ 
    18'h11960: Data = 4'h2; //+ 
    18'h11961: Data = 4'h2; //+ 
    18'h11962: Data = 4'h2; //+ 
    18'h11963: Data = 4'h2; //+ 
    18'h11964: Data = 4'h2; //+ 
    18'h11965: Data = 4'h2; //+ 
    18'h11966: Data = 4'h2; //+ 
    18'h11967: Data = 4'h4; //> 
    18'h11968: Data = 4'h4; //> 
    18'h11969: Data = 4'h6; //[ 
    18'h11970: Data = 4'h3; //- 
    18'h11971: Data = 4'h5; //< 
    18'h11972: Data = 4'h5; //< 
    18'h11973: Data = 4'h5; //< 
    18'h11974: Data = 4'h5; //< 
    18'h11975: Data = 4'h2; //+ 
    18'h11976: Data = 4'h4; //> 
    18'h11977: Data = 4'h4; //> 
    18'h11978: Data = 4'h4; //> 
    18'h11979: Data = 4'h4; //> 
    18'h11980: Data = 4'h7; //] 
    18'h11981: Data = 4'h5; //< 
    18'h11982: Data = 4'h5; //< 
    18'h11983: Data = 4'h5; //< 
    18'h11984: Data = 4'h5; //< 
    18'h11985: Data = 4'h6; //[ 
    18'h11986: Data = 4'h3; //- 
    18'h11987: Data = 4'h4; //> 
    18'h11988: Data = 4'h4; //> 
    18'h11989: Data = 4'h4; //> 
    18'h11990: Data = 4'h4; //> 
    18'h11991: Data = 4'h2; //+ 
    18'h11992: Data = 4'h5; //< 
    18'h11993: Data = 4'h5; //< 
    18'h11994: Data = 4'ha; //0 
    18'h11995: Data = 4'h5; //< 
    18'h11996: Data = 4'h5; //< 
    18'h11997: Data = 4'h7; //] 
    18'h11998: Data = 4'h4; //> 
    18'h11999: Data = 4'h4; //> 
    18'h12000: Data = 4'h6; //[ 
    18'h12001: Data = 4'h5; //< 
    18'h12002: Data = 4'h5; //< 
    18'h12003: Data = 4'h5; //< 
    18'h12004: Data = 4'h5; //< 
    18'h12005: Data = 4'h5; //< 
    18'h12006: Data = 4'h5; //< 
    18'h12007: Data = 4'h5; //< 
    18'h12008: Data = 4'h2; //+ 
    18'h12009: Data = 4'h5; //< 
    18'h12010: Data = 4'h6; //[ 
    18'h12011: Data = 4'h3; //- 
    18'h12012: Data = 4'h5; //< 
    18'h12013: Data = 4'h2; //+ 
    18'h12014: Data = 4'h4; //> 
    18'h12015: Data = 4'h4; //> 
    18'h12016: Data = 4'h4; //> 
    18'h12017: Data = 4'h4; //> 
    18'h12018: Data = 4'h2; //+ 
    18'h12019: Data = 4'h5; //< 
    18'h12020: Data = 4'h5; //< 
    18'h12021: Data = 4'ha; //0 
    18'h12022: Data = 4'h7; //] 
    18'h12023: Data = 4'h4; //> 
    18'h12024: Data = 4'h6; //[ 
    18'h12025: Data = 4'h3; //- 
    18'h12026: Data = 4'h5; //< 
    18'h12027: Data = 4'h5; //< 
    18'h12028: Data = 4'h6; //[ 
    18'h12029: Data = 4'h3; //- 
    18'h12030: Data = 4'h4; //> 
    18'h12031: Data = 4'h2; //+ 
    18'h12032: Data = 4'h4; //> 
    18'h12033: Data = 4'h4; //> 
    18'h12034: Data = 4'h4; //> 
    18'h12035: Data = 4'h3; //- 
    18'h12036: Data = 4'h5; //< 
    18'h12037: Data = 4'h5; //< 
    18'h12038: Data = 4'h5; //< 
    18'h12039: Data = 4'h5; //< 
    18'h12040: Data = 4'h7; //] 
    18'h12041: Data = 4'h4; //> 
    18'h12042: Data = 4'h4; //> 
    18'h12043: Data = 4'h4; //> 
    18'h12044: Data = 4'h7; //] 
    18'h12045: Data = 4'h4; //> 
    18'h12046: Data = 4'h4; //> 
    18'h12047: Data = 4'h4; //> 
    18'h12048: Data = 4'h4; //> 
    18'h12049: Data = 4'h4; //> 
    18'h12050: Data = 4'h4; //> 
    18'h12051: Data = 4'h4; //> 
    18'h12052: Data = 4'h4; //> 
    18'h12053: Data = 4'h4; //> 
    18'h12054: Data = 4'h4; //> 
    18'h12055: Data = 4'h4; //> 
    18'h12056: Data = 4'h4; //> 
    18'h12057: Data = 4'h4; //> 
    18'h12058: Data = 4'h6; //[ 
    18'h12059: Data = 4'h4; //> 
    18'h12060: Data = 4'h4; //> 
    18'h12061: Data = 4'ha; //0 
    18'h12062: Data = 4'h4; //> 
    18'h12063: Data = 4'ha; //0 
    18'h12064: Data = 4'h4; //> 
    18'h12065: Data = 4'ha; //0 
    18'h12066: Data = 4'h4; //> 
    18'h12067: Data = 4'h4; //> 
    18'h12068: Data = 4'h4; //> 
    18'h12069: Data = 4'h4; //> 
    18'h12070: Data = 4'h4; //> 
    18'h12071: Data = 4'h7; //] 
    18'h12072: Data = 4'h5; //< 
    18'h12073: Data = 4'h5; //< 
    18'h12074: Data = 4'h5; //< 
    18'h12075: Data = 4'h5; //< 
    18'h12076: Data = 4'h5; //< 
    18'h12077: Data = 4'h5; //< 
    18'h12078: Data = 4'h5; //< 
    18'h12079: Data = 4'h5; //< 
    18'h12080: Data = 4'h5; //< 
    18'h12081: Data = 4'h6; //[ 
    18'h12082: Data = 4'h5; //< 
    18'h12083: Data = 4'h5; //< 
    18'h12084: Data = 4'h5; //< 
    18'h12085: Data = 4'h5; //< 
    18'h12086: Data = 4'h5; //< 
    18'h12087: Data = 4'h5; //< 
    18'h12088: Data = 4'h5; //< 
    18'h12089: Data = 4'h5; //< 
    18'h12090: Data = 4'h5; //< 
    18'h12091: Data = 4'h7; //] 
    18'h12092: Data = 4'h4; //> 
    18'h12093: Data = 4'h4; //> 
    18'h12094: Data = 4'h4; //> 
    18'h12095: Data = 4'ha; //0 
    18'h12096: Data = 4'h4; //> 
    18'h12097: Data = 4'h4; //> 
    18'h12098: Data = 4'h4; //> 
    18'h12099: Data = 4'h4; //> 
    18'h12100: Data = 4'h4; //> 
    18'h12101: Data = 4'h4; //> 
    18'h12102: Data = 4'h6; //[ 
    18'h12103: Data = 4'h4; //> 
    18'h12104: Data = 4'h4; //> 
    18'h12105: Data = 4'h4; //> 
    18'h12106: Data = 4'h4; //> 
    18'h12107: Data = 4'h4; //> 
    18'h12108: Data = 4'h6; //[ 
    18'h12109: Data = 4'h3; //- 
    18'h12110: Data = 4'h5; //< 
    18'h12111: Data = 4'h5; //< 
    18'h12112: Data = 4'h5; //< 
    18'h12113: Data = 4'h5; //< 
    18'h12114: Data = 4'h2; //+ 
    18'h12115: Data = 4'h4; //> 
    18'h12116: Data = 4'h4; //> 
    18'h12117: Data = 4'h4; //> 
    18'h12118: Data = 4'h4; //> 
    18'h12119: Data = 4'h7; //] 
    18'h12120: Data = 4'h5; //< 
    18'h12121: Data = 4'h5; //< 
    18'h12122: Data = 4'h5; //< 
    18'h12123: Data = 4'h5; //< 
    18'h12124: Data = 4'h6; //[ 
    18'h12125: Data = 4'h3; //- 
    18'h12126: Data = 4'h4; //> 
    18'h12127: Data = 4'h4; //> 
    18'h12128: Data = 4'h4; //> 
    18'h12129: Data = 4'h4; //> 
    18'h12130: Data = 4'h2; //+ 
    18'h12131: Data = 4'h5; //< 
    18'h12132: Data = 4'h5; //< 
    18'h12133: Data = 4'h5; //< 
    18'h12134: Data = 4'h2; //+ 
    18'h12135: Data = 4'h5; //< 
    18'h12136: Data = 4'h7; //] 
    18'h12137: Data = 4'h4; //> 
    18'h12138: Data = 4'h4; //> 
    18'h12139: Data = 4'h4; //> 
    18'h12140: Data = 4'h4; //> 
    18'h12141: Data = 4'h4; //> 
    18'h12142: Data = 4'h4; //> 
    18'h12143: Data = 4'h4; //> 
    18'h12144: Data = 4'h4; //> 
    18'h12145: Data = 4'h7; //] 
    18'h12146: Data = 4'h5; //< 
    18'h12147: Data = 4'h5; //< 
    18'h12148: Data = 4'h5; //< 
    18'h12149: Data = 4'h5; //< 
    18'h12150: Data = 4'h5; //< 
    18'h12151: Data = 4'h5; //< 
    18'h12152: Data = 4'h5; //< 
    18'h12153: Data = 4'h5; //< 
    18'h12154: Data = 4'h5; //< 
    18'h12155: Data = 4'h6; //[ 
    18'h12156: Data = 4'h5; //< 
    18'h12157: Data = 4'h5; //< 
    18'h12158: Data = 4'h5; //< 
    18'h12159: Data = 4'h5; //< 
    18'h12160: Data = 4'h5; //< 
    18'h12161: Data = 4'h5; //< 
    18'h12162: Data = 4'h5; //< 
    18'h12163: Data = 4'h5; //< 
    18'h12164: Data = 4'h5; //< 
    18'h12165: Data = 4'h7; //] 
    18'h12166: Data = 4'h4; //> 
    18'h12167: Data = 4'h4; //> 
    18'h12168: Data = 4'h4; //> 
    18'h12169: Data = 4'h4; //> 
    18'h12170: Data = 4'h4; //> 
    18'h12171: Data = 4'h4; //> 
    18'h12172: Data = 4'h4; //> 
    18'h12173: Data = 4'h4; //> 
    18'h12174: Data = 4'h4; //> 
    18'h12175: Data = 4'h6; //[ 
    18'h12176: Data = 4'h4; //> 
    18'h12177: Data = 4'h4; //> 
    18'h12178: Data = 4'h6; //[ 
    18'h12179: Data = 4'h3; //- 
    18'h12180: Data = 4'h5; //< 
    18'h12181: Data = 4'h5; //< 
    18'h12182: Data = 4'h5; //< 
    18'h12183: Data = 4'h5; //< 
    18'h12184: Data = 4'h5; //< 
    18'h12185: Data = 4'h5; //< 
    18'h12186: Data = 4'h5; //< 
    18'h12187: Data = 4'h5; //< 
    18'h12188: Data = 4'h5; //< 
    18'h12189: Data = 4'h2; //+ 
    18'h12190: Data = 4'h4; //> 
    18'h12191: Data = 4'h4; //> 
    18'h12192: Data = 4'h4; //> 
    18'h12193: Data = 4'h4; //> 
    18'h12194: Data = 4'h4; //> 
    18'h12195: Data = 4'h4; //> 
    18'h12196: Data = 4'h4; //> 
    18'h12197: Data = 4'h4; //> 
    18'h12198: Data = 4'h4; //> 
    18'h12199: Data = 4'h7; //] 
    18'h12200: Data = 4'h4; //> 
    18'h12201: Data = 4'h4; //> 
    18'h12202: Data = 4'h4; //> 
    18'h12203: Data = 4'h4; //> 
    18'h12204: Data = 4'h4; //> 
    18'h12205: Data = 4'h4; //> 
    18'h12206: Data = 4'h4; //> 
    18'h12207: Data = 4'h7; //] 
    18'h12208: Data = 4'h5; //< 
    18'h12209: Data = 4'h5; //< 
    18'h12210: Data = 4'h5; //< 
    18'h12211: Data = 4'h5; //< 
    18'h12212: Data = 4'h5; //< 
    18'h12213: Data = 4'h5; //< 
    18'h12214: Data = 4'h5; //< 
    18'h12215: Data = 4'h5; //< 
    18'h12216: Data = 4'h5; //< 
    18'h12217: Data = 4'h6; //[ 
    18'h12218: Data = 4'h5; //< 
    18'h12219: Data = 4'h5; //< 
    18'h12220: Data = 4'h5; //< 
    18'h12221: Data = 4'h5; //< 
    18'h12222: Data = 4'h5; //< 
    18'h12223: Data = 4'h5; //< 
    18'h12224: Data = 4'h5; //< 
    18'h12225: Data = 4'h5; //< 
    18'h12226: Data = 4'h5; //< 
    18'h12227: Data = 4'h7; //] 
    18'h12228: Data = 4'h4; //> 
    18'h12229: Data = 4'h4; //> 
    18'h12230: Data = 4'h4; //> 
    18'h12231: Data = 4'h4; //> 
    18'h12232: Data = 4'h4; //> 
    18'h12233: Data = 4'h4; //> 
    18'h12234: Data = 4'h4; //> 
    18'h12235: Data = 4'h4; //> 
    18'h12236: Data = 4'h4; //> 
    18'h12237: Data = 4'h2; //+ 
    18'h12238: Data = 4'h2; //+ 
    18'h12239: Data = 4'h2; //+ 
    18'h12240: Data = 4'h2; //+ 
    18'h12241: Data = 4'h2; //+ 
    18'h12242: Data = 4'h2; //+ 
    18'h12243: Data = 4'h2; //+ 
    18'h12244: Data = 4'h2; //+ 
    18'h12245: Data = 4'h2; //+ 
    18'h12246: Data = 4'h2; //+ 
    18'h12247: Data = 4'h2; //+ 
    18'h12248: Data = 4'h2; //+ 
    18'h12249: Data = 4'h2; //+ 
    18'h12250: Data = 4'h2; //+ 
    18'h12251: Data = 4'h2; //+ 
    18'h12252: Data = 4'h6; //[ 
    18'h12253: Data = 4'h6; //[ 
    18'h12254: Data = 4'h4; //> 
    18'h12255: Data = 4'h4; //> 
    18'h12256: Data = 4'h4; //> 
    18'h12257: Data = 4'h4; //> 
    18'h12258: Data = 4'h4; //> 
    18'h12259: Data = 4'h4; //> 
    18'h12260: Data = 4'h4; //> 
    18'h12261: Data = 4'h4; //> 
    18'h12262: Data = 4'h4; //> 
    18'h12263: Data = 4'h7; //] 
    18'h12264: Data = 4'h2; //+ 
    18'h12265: Data = 4'h4; //> 
    18'h12266: Data = 4'h6; //[ 
    18'h12267: Data = 4'h3; //- 
    18'h12268: Data = 4'h7; //] 
    18'h12269: Data = 4'h4; //> 
    18'h12270: Data = 4'ha; //0 
    18'h12271: Data = 4'h4; //> 
    18'h12272: Data = 4'ha; //0 
    18'h12273: Data = 4'h4; //> 
    18'h12274: Data = 4'ha; //0 
    18'h12275: Data = 4'h4; //> 
    18'h12276: Data = 4'ha; //0 
    18'h12277: Data = 4'h4; //> 
    18'h12278: Data = 4'ha; //0 
    18'h12279: Data = 4'h4; //> 
    18'h12280: Data = 4'ha; //0 
    18'h12281: Data = 4'h4; //> 
    18'h12282: Data = 4'ha; //0 
    18'h12283: Data = 4'h4; //> 
    18'h12284: Data = 4'ha; //0 
    18'h12285: Data = 4'h5; //< 
    18'h12286: Data = 4'h5; //< 
    18'h12287: Data = 4'h5; //< 
    18'h12288: Data = 4'h5; //< 
    18'h12289: Data = 4'h5; //< 
    18'h12290: Data = 4'h5; //< 
    18'h12291: Data = 4'h5; //< 
    18'h12292: Data = 4'h5; //< 
    18'h12293: Data = 4'h5; //< 
    18'h12294: Data = 4'h6; //[ 
    18'h12295: Data = 4'h5; //< 
    18'h12296: Data = 4'h5; //< 
    18'h12297: Data = 4'h5; //< 
    18'h12298: Data = 4'h5; //< 
    18'h12299: Data = 4'h5; //< 
    18'h12300: Data = 4'h5; //< 
    18'h12301: Data = 4'h5; //< 
    18'h12302: Data = 4'h5; //< 
    18'h12303: Data = 4'h5; //< 
    18'h12304: Data = 4'h7; //] 
    18'h12305: Data = 4'h4; //> 
    18'h12306: Data = 4'h4; //> 
    18'h12307: Data = 4'h4; //> 
    18'h12308: Data = 4'h4; //> 
    18'h12309: Data = 4'h4; //> 
    18'h12310: Data = 4'h4; //> 
    18'h12311: Data = 4'h4; //> 
    18'h12312: Data = 4'h4; //> 
    18'h12313: Data = 4'h4; //> 
    18'h12314: Data = 4'h3; //- 
    18'h12315: Data = 4'h7; //] 
    18'h12316: Data = 4'h2; //+ 
    18'h12317: Data = 4'h6; //[ 
    18'h12318: Data = 4'h4; //> 
    18'h12319: Data = 4'h2; //+ 
    18'h12320: Data = 4'h4; //> 
    18'h12321: Data = 4'h4; //> 
    18'h12322: Data = 4'h4; //> 
    18'h12323: Data = 4'h4; //> 
    18'h12324: Data = 4'h4; //> 
    18'h12325: Data = 4'h4; //> 
    18'h12326: Data = 4'h4; //> 
    18'h12327: Data = 4'h4; //> 
    18'h12328: Data = 4'h7; //] 
    18'h12329: Data = 4'h5; //< 
    18'h12330: Data = 4'h5; //< 
    18'h12331: Data = 4'h5; //< 
    18'h12332: Data = 4'h5; //< 
    18'h12333: Data = 4'h5; //< 
    18'h12334: Data = 4'h5; //< 
    18'h12335: Data = 4'h5; //< 
    18'h12336: Data = 4'h5; //< 
    18'h12337: Data = 4'h5; //< 
    18'h12338: Data = 4'h6; //[ 
    18'h12339: Data = 4'h5; //< 
    18'h12340: Data = 4'h5; //< 
    18'h12341: Data = 4'h5; //< 
    18'h12342: Data = 4'h5; //< 
    18'h12343: Data = 4'h5; //< 
    18'h12344: Data = 4'h5; //< 
    18'h12345: Data = 4'h5; //< 
    18'h12346: Data = 4'h5; //< 
    18'h12347: Data = 4'h5; //< 
    18'h12348: Data = 4'h7; //] 
    18'h12349: Data = 4'h4; //> 
    18'h12350: Data = 4'h4; //> 
    18'h12351: Data = 4'h4; //> 
    18'h12352: Data = 4'h4; //> 
    18'h12353: Data = 4'h4; //> 
    18'h12354: Data = 4'h4; //> 
    18'h12355: Data = 4'h4; //> 
    18'h12356: Data = 4'h4; //> 
    18'h12357: Data = 4'h4; //> 
    18'h12358: Data = 4'h6; //[ 
    18'h12359: Data = 4'h4; //> 
    18'h12360: Data = 4'h3; //- 
    18'h12361: Data = 4'h4; //> 
    18'h12362: Data = 4'h4; //> 
    18'h12363: Data = 4'h4; //> 
    18'h12364: Data = 4'h4; //> 
    18'h12365: Data = 4'h4; //> 
    18'h12366: Data = 4'h6; //[ 
    18'h12367: Data = 4'h3; //- 
    18'h12368: Data = 4'h5; //< 
    18'h12369: Data = 4'h5; //< 
    18'h12370: Data = 4'h5; //< 
    18'h12371: Data = 4'h5; //< 
    18'h12372: Data = 4'h5; //< 
    18'h12373: Data = 4'h2; //+ 
    18'h12374: Data = 4'h4; //> 
    18'h12375: Data = 4'h4; //> 
    18'h12376: Data = 4'h4; //> 
    18'h12377: Data = 4'h4; //> 
    18'h12378: Data = 4'h4; //> 
    18'h12379: Data = 4'h7; //] 
    18'h12380: Data = 4'h5; //< 
    18'h12381: Data = 4'h5; //< 
    18'h12382: Data = 4'h5; //< 
    18'h12383: Data = 4'h5; //< 
    18'h12384: Data = 4'h5; //< 
    18'h12385: Data = 4'h6; //[ 
    18'h12386: Data = 4'h3; //- 
    18'h12387: Data = 4'h4; //> 
    18'h12388: Data = 4'h4; //> 
    18'h12389: Data = 4'h4; //> 
    18'h12390: Data = 4'h4; //> 
    18'h12391: Data = 4'h4; //> 
    18'h12392: Data = 4'h2; //+ 
    18'h12393: Data = 4'h5; //< 
    18'h12394: Data = 4'h5; //< 
    18'h12395: Data = 4'h5; //< 
    18'h12396: Data = 4'h5; //< 
    18'h12397: Data = 4'h5; //< 
    18'h12398: Data = 4'h5; //< 
    18'h12399: Data = 4'h6; //[ 
    18'h12400: Data = 4'h3; //- 
    18'h12401: Data = 4'h4; //> 
    18'h12402: Data = 4'h4; //> 
    18'h12403: Data = 4'h6; //[ 
    18'h12404: Data = 4'h3; //- 
    18'h12405: Data = 4'h5; //< 
    18'h12406: Data = 4'h5; //< 
    18'h12407: Data = 4'h2; //+ 
    18'h12408: Data = 4'h4; //> 
    18'h12409: Data = 4'h4; //> 
    18'h12410: Data = 4'h7; //] 
    18'h12411: Data = 4'h5; //< 
    18'h12412: Data = 4'h5; //< 
    18'h12413: Data = 4'h6; //[ 
    18'h12414: Data = 4'h3; //- 
    18'h12415: Data = 4'h4; //> 
    18'h12416: Data = 4'h4; //> 
    18'h12417: Data = 4'h2; //+ 
    18'h12418: Data = 4'h4; //> 
    18'h12419: Data = 4'h2; //+ 
    18'h12420: Data = 4'h5; //< 
    18'h12421: Data = 4'h5; //< 
    18'h12422: Data = 4'h5; //< 
    18'h12423: Data = 4'h7; //] 
    18'h12424: Data = 4'h2; //+ 
    18'h12425: Data = 4'h4; //> 
    18'h12426: Data = 4'h4; //> 
    18'h12427: Data = 4'h4; //> 
    18'h12428: Data = 4'h4; //> 
    18'h12429: Data = 4'h4; //> 
    18'h12430: Data = 4'h4; //> 
    18'h12431: Data = 4'h4; //> 
    18'h12432: Data = 4'h4; //> 
    18'h12433: Data = 4'h4; //> 
    18'h12434: Data = 4'h7; //] 
    18'h12435: Data = 4'h5; //< 
    18'h12436: Data = 4'h5; //< 
    18'h12437: Data = 4'h5; //< 
    18'h12438: Data = 4'h5; //< 
    18'h12439: Data = 4'h5; //< 
    18'h12440: Data = 4'h5; //< 
    18'h12441: Data = 4'h5; //< 
    18'h12442: Data = 4'h5; //< 
    18'h12443: Data = 4'h6; //[ 
    18'h12444: Data = 4'h5; //< 
    18'h12445: Data = 4'h5; //< 
    18'h12446: Data = 4'h5; //< 
    18'h12447: Data = 4'h5; //< 
    18'h12448: Data = 4'h5; //< 
    18'h12449: Data = 4'h5; //< 
    18'h12450: Data = 4'h5; //< 
    18'h12451: Data = 4'h5; //< 
    18'h12452: Data = 4'h5; //< 
    18'h12453: Data = 4'h7; //] 
    18'h12454: Data = 4'h7; //] 
    18'h12455: Data = 4'h4; //> 
    18'h12456: Data = 4'h4; //> 
    18'h12457: Data = 4'h4; //> 
    18'h12458: Data = 4'h4; //> 
    18'h12459: Data = 4'h4; //> 
    18'h12460: Data = 4'h4; //> 
    18'h12461: Data = 4'h4; //> 
    18'h12462: Data = 4'h4; //> 
    18'h12463: Data = 4'h4; //> 
    18'h12464: Data = 4'h6; //[ 
    18'h12465: Data = 4'h4; //> 
    18'h12466: Data = 4'h4; //> 
    18'h12467: Data = 4'h4; //> 
    18'h12468: Data = 4'h4; //> 
    18'h12469: Data = 4'h4; //> 
    18'h12470: Data = 4'h4; //> 
    18'h12471: Data = 4'h4; //> 
    18'h12472: Data = 4'h4; //> 
    18'h12473: Data = 4'h4; //> 
    18'h12474: Data = 4'h7; //] 
    18'h12475: Data = 4'h5; //< 
    18'h12476: Data = 4'h5; //< 
    18'h12477: Data = 4'h5; //< 
    18'h12478: Data = 4'h5; //< 
    18'h12479: Data = 4'h5; //< 
    18'h12480: Data = 4'h5; //< 
    18'h12481: Data = 4'h5; //< 
    18'h12482: Data = 4'h5; //< 
    18'h12483: Data = 4'h5; //< 
    18'h12484: Data = 4'h6; //[ 
    18'h12485: Data = 4'h4; //> 
    18'h12486: Data = 4'h6; //[ 
    18'h12487: Data = 4'h3; //- 
    18'h12488: Data = 4'h4; //> 
    18'h12489: Data = 4'h4; //> 
    18'h12490: Data = 4'h4; //> 
    18'h12491: Data = 4'h4; //> 
    18'h12492: Data = 4'h4; //> 
    18'h12493: Data = 4'h4; //> 
    18'h12494: Data = 4'h4; //> 
    18'h12495: Data = 4'h4; //> 
    18'h12496: Data = 4'h4; //> 
    18'h12497: Data = 4'h2; //+ 
    18'h12498: Data = 4'h5; //< 
    18'h12499: Data = 4'h5; //< 
    18'h12500: Data = 4'h5; //< 
    18'h12501: Data = 4'h5; //< 
    18'h12502: Data = 4'h5; //< 
    18'h12503: Data = 4'h5; //< 
    18'h12504: Data = 4'h5; //< 
    18'h12505: Data = 4'h5; //< 
    18'h12506: Data = 4'h5; //< 
    18'h12507: Data = 4'h7; //] 
    18'h12508: Data = 4'h5; //< 
    18'h12509: Data = 4'h5; //< 
    18'h12510: Data = 4'h5; //< 
    18'h12511: Data = 4'h5; //< 
    18'h12512: Data = 4'h5; //< 
    18'h12513: Data = 4'h5; //< 
    18'h12514: Data = 4'h5; //< 
    18'h12515: Data = 4'h5; //< 
    18'h12516: Data = 4'h5; //< 
    18'h12517: Data = 4'h5; //< 
    18'h12518: Data = 4'h7; //] 
    18'h12519: Data = 4'h4; //> 
    18'h12520: Data = 4'h6; //[ 
    18'h12521: Data = 4'h3; //- 
    18'h12522: Data = 4'h4; //> 
    18'h12523: Data = 4'h4; //> 
    18'h12524: Data = 4'h4; //> 
    18'h12525: Data = 4'h4; //> 
    18'h12526: Data = 4'h4; //> 
    18'h12527: Data = 4'h4; //> 
    18'h12528: Data = 4'h4; //> 
    18'h12529: Data = 4'h4; //> 
    18'h12530: Data = 4'h4; //> 
    18'h12531: Data = 4'h2; //+ 
    18'h12532: Data = 4'h5; //< 
    18'h12533: Data = 4'h5; //< 
    18'h12534: Data = 4'h5; //< 
    18'h12535: Data = 4'h5; //< 
    18'h12536: Data = 4'h5; //< 
    18'h12537: Data = 4'h5; //< 
    18'h12538: Data = 4'h5; //< 
    18'h12539: Data = 4'h5; //< 
    18'h12540: Data = 4'h5; //< 
    18'h12541: Data = 4'h7; //] 
    18'h12542: Data = 4'h5; //< 
    18'h12543: Data = 4'h2; //+ 
    18'h12544: Data = 4'h4; //> 
    18'h12545: Data = 4'h4; //> 
    18'h12546: Data = 4'h4; //> 
    18'h12547: Data = 4'h4; //> 
    18'h12548: Data = 4'h4; //> 
    18'h12549: Data = 4'h4; //> 
    18'h12550: Data = 4'h4; //> 
    18'h12551: Data = 4'h4; //> 
    18'h12552: Data = 4'h7; //] 
    18'h12553: Data = 4'h5; //< 
    18'h12554: Data = 4'h5; //< 
    18'h12555: Data = 4'h5; //< 
    18'h12556: Data = 4'h5; //< 
    18'h12557: Data = 4'h5; //< 
    18'h12558: Data = 4'h5; //< 
    18'h12559: Data = 4'h5; //< 
    18'h12560: Data = 4'h5; //< 
    18'h12561: Data = 4'h5; //< 
    18'h12562: Data = 4'h6; //[ 
    18'h12563: Data = 4'h4; //> 
    18'h12564: Data = 4'ha; //0 
    18'h12565: Data = 4'h5; //< 
    18'h12566: Data = 4'h3; //- 
    18'h12567: Data = 4'h4; //> 
    18'h12568: Data = 4'h4; //> 
    18'h12569: Data = 4'h4; //> 
    18'h12570: Data = 4'h6; //[ 
    18'h12571: Data = 4'h3; //- 
    18'h12572: Data = 4'h5; //< 
    18'h12573: Data = 4'h5; //< 
    18'h12574: Data = 4'h5; //< 
    18'h12575: Data = 4'h2; //+ 
    18'h12576: Data = 4'h4; //> 
    18'h12577: Data = 4'h6; //[ 
    18'h12578: Data = 4'h5; //< 
    18'h12579: Data = 4'h3; //- 
    18'h12580: Data = 4'h4; //> 
    18'h12581: Data = 4'h3; //- 
    18'h12582: Data = 4'h5; //< 
    18'h12583: Data = 4'h5; //< 
    18'h12584: Data = 4'h5; //< 
    18'h12585: Data = 4'h5; //< 
    18'h12586: Data = 4'h5; //< 
    18'h12587: Data = 4'h5; //< 
    18'h12588: Data = 4'h5; //< 
    18'h12589: Data = 4'h2; //+ 
    18'h12590: Data = 4'h4; //> 
    18'h12591: Data = 4'h4; //> 
    18'h12592: Data = 4'h4; //> 
    18'h12593: Data = 4'h4; //> 
    18'h12594: Data = 4'h4; //> 
    18'h12595: Data = 4'h4; //> 
    18'h12596: Data = 4'h4; //> 
    18'h12597: Data = 4'h7; //] 
    18'h12598: Data = 4'h5; //< 
    18'h12599: Data = 4'h6; //[ 
    18'h12600: Data = 4'h3; //- 
    18'h12601: Data = 4'h4; //> 
    18'h12602: Data = 4'h2; //+ 
    18'h12603: Data = 4'h5; //< 
    18'h12604: Data = 4'h7; //] 
    18'h12605: Data = 4'h4; //> 
    18'h12606: Data = 4'h4; //> 
    18'h12607: Data = 4'h4; //> 
    18'h12608: Data = 4'h7; //] 
    18'h12609: Data = 4'h5; //< 
    18'h12610: Data = 4'h5; //< 
    18'h12611: Data = 4'h6; //[ 
    18'h12612: Data = 4'h3; //- 
    18'h12613: Data = 4'h4; //> 
    18'h12614: Data = 4'h4; //> 
    18'h12615: Data = 4'h2; //+ 
    18'h12616: Data = 4'h5; //< 
    18'h12617: Data = 4'h5; //< 
    18'h12618: Data = 4'h7; //] 
    18'h12619: Data = 4'h5; //< 
    18'h12620: Data = 4'h2; //+ 
    18'h12621: Data = 4'h5; //< 
    18'h12622: Data = 4'h5; //< 
    18'h12623: Data = 4'h5; //< 
    18'h12624: Data = 4'h5; //< 
    18'h12625: Data = 4'h5; //< 
    18'h12626: Data = 4'h5; //< 
    18'h12627: Data = 4'h5; //< 
    18'h12628: Data = 4'h5; //< 
    18'h12629: Data = 4'h5; //< 
    18'h12630: Data = 4'h7; //] 
    18'h12631: Data = 4'h4; //> 
    18'h12632: Data = 4'h4; //> 
    18'h12633: Data = 4'h4; //> 
    18'h12634: Data = 4'h4; //> 
    18'h12635: Data = 4'h4; //> 
    18'h12636: Data = 4'h4; //> 
    18'h12637: Data = 4'h4; //> 
    18'h12638: Data = 4'h4; //> 
    18'h12639: Data = 4'h4; //> 
    18'h12640: Data = 4'h6; //[ 
    18'h12641: Data = 4'h4; //> 
    18'h12642: Data = 4'h4; //> 
    18'h12643: Data = 4'h4; //> 
    18'h12644: Data = 4'h4; //> 
    18'h12645: Data = 4'h4; //> 
    18'h12646: Data = 4'h4; //> 
    18'h12647: Data = 4'h6; //[ 
    18'h12648: Data = 4'h3; //- 
    18'h12649: Data = 4'h5; //< 
    18'h12650: Data = 4'h5; //< 
    18'h12651: Data = 4'h5; //< 
    18'h12652: Data = 4'h5; //< 
    18'h12653: Data = 4'h5; //< 
    18'h12654: Data = 4'h2; //+ 
    18'h12655: Data = 4'h4; //> 
    18'h12656: Data = 4'h4; //> 
    18'h12657: Data = 4'h4; //> 
    18'h12658: Data = 4'h4; //> 
    18'h12659: Data = 4'h4; //> 
    18'h12660: Data = 4'h7; //] 
    18'h12661: Data = 4'h5; //< 
    18'h12662: Data = 4'h5; //< 
    18'h12663: Data = 4'h5; //< 
    18'h12664: Data = 4'h5; //< 
    18'h12665: Data = 4'h5; //< 
    18'h12666: Data = 4'h6; //[ 
    18'h12667: Data = 4'h3; //- 
    18'h12668: Data = 4'h4; //> 
    18'h12669: Data = 4'h4; //> 
    18'h12670: Data = 4'h4; //> 
    18'h12671: Data = 4'h4; //> 
    18'h12672: Data = 4'h4; //> 
    18'h12673: Data = 4'h2; //+ 
    18'h12674: Data = 4'h5; //< 
    18'h12675: Data = 4'h5; //< 
    18'h12676: Data = 4'h5; //< 
    18'h12677: Data = 4'h5; //< 
    18'h12678: Data = 4'h2; //+ 
    18'h12679: Data = 4'h5; //< 
    18'h12680: Data = 4'h7; //] 
    18'h12681: Data = 4'h4; //> 
    18'h12682: Data = 4'h4; //> 
    18'h12683: Data = 4'h4; //> 
    18'h12684: Data = 4'h4; //> 
    18'h12685: Data = 4'h4; //> 
    18'h12686: Data = 4'h4; //> 
    18'h12687: Data = 4'h4; //> 
    18'h12688: Data = 4'h4; //> 
    18'h12689: Data = 4'h7; //] 
    18'h12690: Data = 4'h5; //< 
    18'h12691: Data = 4'h5; //< 
    18'h12692: Data = 4'h5; //< 
    18'h12693: Data = 4'h5; //< 
    18'h12694: Data = 4'h5; //< 
    18'h12695: Data = 4'h5; //< 
    18'h12696: Data = 4'h5; //< 
    18'h12697: Data = 4'h5; //< 
    18'h12698: Data = 4'h5; //< 
    18'h12699: Data = 4'h6; //[ 
    18'h12700: Data = 4'h5; //< 
    18'h12701: Data = 4'h5; //< 
    18'h12702: Data = 4'h5; //< 
    18'h12703: Data = 4'h5; //< 
    18'h12704: Data = 4'h5; //< 
    18'h12705: Data = 4'h5; //< 
    18'h12706: Data = 4'h5; //< 
    18'h12707: Data = 4'h5; //< 
    18'h12708: Data = 4'h5; //< 
    18'h12709: Data = 4'h7; //] 
    18'h12710: Data = 4'h4; //> 
    18'h12711: Data = 4'h4; //> 
    18'h12712: Data = 4'h4; //> 
    18'h12713: Data = 4'h4; //> 
    18'h12714: Data = 4'h4; //> 
    18'h12715: Data = 4'h4; //> 
    18'h12716: Data = 4'h4; //> 
    18'h12717: Data = 4'h4; //> 
    18'h12718: Data = 4'h4; //> 
    18'h12719: Data = 4'h6; //[ 
    18'h12720: Data = 4'h4; //> 
    18'h12721: Data = 4'h2; //+ 
    18'h12722: Data = 4'h4; //> 
    18'h12723: Data = 4'h4; //> 
    18'h12724: Data = 4'h4; //> 
    18'h12725: Data = 4'h4; //> 
    18'h12726: Data = 4'h4; //> 
    18'h12727: Data = 4'h4; //> 
    18'h12728: Data = 4'h4; //> 
    18'h12729: Data = 4'h4; //> 
    18'h12730: Data = 4'h7; //] 
    18'h12731: Data = 4'h5; //< 
    18'h12732: Data = 4'h5; //< 
    18'h12733: Data = 4'h5; //< 
    18'h12734: Data = 4'h5; //< 
    18'h12735: Data = 4'h5; //< 
    18'h12736: Data = 4'h5; //< 
    18'h12737: Data = 4'h5; //< 
    18'h12738: Data = 4'h5; //< 
    18'h12739: Data = 4'h5; //< 
    18'h12740: Data = 4'h6; //[ 
    18'h12741: Data = 4'h5; //< 
    18'h12742: Data = 4'h5; //< 
    18'h12743: Data = 4'h5; //< 
    18'h12744: Data = 4'h5; //< 
    18'h12745: Data = 4'h5; //< 
    18'h12746: Data = 4'h5; //< 
    18'h12747: Data = 4'h5; //< 
    18'h12748: Data = 4'h5; //< 
    18'h12749: Data = 4'h5; //< 
    18'h12750: Data = 4'h7; //] 
    18'h12751: Data = 4'h4; //> 
    18'h12752: Data = 4'h4; //> 
    18'h12753: Data = 4'h4; //> 
    18'h12754: Data = 4'h4; //> 
    18'h12755: Data = 4'h4; //> 
    18'h12756: Data = 4'h4; //> 
    18'h12757: Data = 4'h4; //> 
    18'h12758: Data = 4'h4; //> 
    18'h12759: Data = 4'h4; //> 
    18'h12760: Data = 4'h6; //[ 
    18'h12761: Data = 4'h4; //> 
    18'h12762: Data = 4'h3; //- 
    18'h12763: Data = 4'h4; //> 
    18'h12764: Data = 4'h4; //> 
    18'h12765: Data = 4'h4; //> 
    18'h12766: Data = 4'h4; //> 
    18'h12767: Data = 4'h4; //> 
    18'h12768: Data = 4'h6; //[ 
    18'h12769: Data = 4'h3; //- 
    18'h12770: Data = 4'h5; //< 
    18'h12771: Data = 4'h5; //< 
    18'h12772: Data = 4'h5; //< 
    18'h12773: Data = 4'h5; //< 
    18'h12774: Data = 4'h5; //< 
    18'h12775: Data = 4'h2; //+ 
    18'h12776: Data = 4'h4; //> 
    18'h12777: Data = 4'h4; //> 
    18'h12778: Data = 4'h4; //> 
    18'h12779: Data = 4'h4; //> 
    18'h12780: Data = 4'h4; //> 
    18'h12781: Data = 4'h7; //] 
    18'h12782: Data = 4'h5; //< 
    18'h12783: Data = 4'h5; //< 
    18'h12784: Data = 4'h5; //< 
    18'h12785: Data = 4'h5; //< 
    18'h12786: Data = 4'h5; //< 
    18'h12787: Data = 4'h6; //[ 
    18'h12788: Data = 4'h3; //- 
    18'h12789: Data = 4'h4; //> 
    18'h12790: Data = 4'h4; //> 
    18'h12791: Data = 4'h4; //> 
    18'h12792: Data = 4'h4; //> 
    18'h12793: Data = 4'h4; //> 
    18'h12794: Data = 4'h2; //+ 
    18'h12795: Data = 4'h5; //< 
    18'h12796: Data = 4'h5; //< 
    18'h12797: Data = 4'h5; //< 
    18'h12798: Data = 4'h5; //< 
    18'h12799: Data = 4'h5; //< 
    18'h12800: Data = 4'h5; //< 
    18'h12801: Data = 4'h6; //[ 
    18'h12802: Data = 4'h3; //- 
    18'h12803: Data = 4'h4; //> 
    18'h12804: Data = 4'h4; //> 
    18'h12805: Data = 4'h6; //[ 
    18'h12806: Data = 4'h3; //- 
    18'h12807: Data = 4'h5; //< 
    18'h12808: Data = 4'h5; //< 
    18'h12809: Data = 4'h2; //+ 
    18'h12810: Data = 4'h4; //> 
    18'h12811: Data = 4'h4; //> 
    18'h12812: Data = 4'h7; //] 
    18'h12813: Data = 4'h5; //< 
    18'h12814: Data = 4'h5; //< 
    18'h12815: Data = 4'h6; //[ 
    18'h12816: Data = 4'h3; //- 
    18'h12817: Data = 4'h4; //> 
    18'h12818: Data = 4'h4; //> 
    18'h12819: Data = 4'h2; //+ 
    18'h12820: Data = 4'h4; //> 
    18'h12821: Data = 4'h4; //> 
    18'h12822: Data = 4'h2; //+ 
    18'h12823: Data = 4'h5; //< 
    18'h12824: Data = 4'h5; //< 
    18'h12825: Data = 4'h5; //< 
    18'h12826: Data = 4'h5; //< 
    18'h12827: Data = 4'h7; //] 
    18'h12828: Data = 4'h2; //+ 
    18'h12829: Data = 4'h4; //> 
    18'h12830: Data = 4'h4; //> 
    18'h12831: Data = 4'h4; //> 
    18'h12832: Data = 4'h4; //> 
    18'h12833: Data = 4'h4; //> 
    18'h12834: Data = 4'h4; //> 
    18'h12835: Data = 4'h4; //> 
    18'h12836: Data = 4'h4; //> 
    18'h12837: Data = 4'h4; //> 
    18'h12838: Data = 4'h7; //] 
    18'h12839: Data = 4'h5; //< 
    18'h12840: Data = 4'h5; //< 
    18'h12841: Data = 4'h5; //< 
    18'h12842: Data = 4'h5; //< 
    18'h12843: Data = 4'h5; //< 
    18'h12844: Data = 4'h5; //< 
    18'h12845: Data = 4'h5; //< 
    18'h12846: Data = 4'h5; //< 
    18'h12847: Data = 4'h6; //[ 
    18'h12848: Data = 4'h5; //< 
    18'h12849: Data = 4'h5; //< 
    18'h12850: Data = 4'h5; //< 
    18'h12851: Data = 4'h5; //< 
    18'h12852: Data = 4'h5; //< 
    18'h12853: Data = 4'h5; //< 
    18'h12854: Data = 4'h5; //< 
    18'h12855: Data = 4'h5; //< 
    18'h12856: Data = 4'h5; //< 
    18'h12857: Data = 4'h7; //] 
    18'h12858: Data = 4'h7; //] 
    18'h12859: Data = 4'h4; //> 
    18'h12860: Data = 4'h4; //> 
    18'h12861: Data = 4'h4; //> 
    18'h12862: Data = 4'h4; //> 
    18'h12863: Data = 4'h4; //> 
    18'h12864: Data = 4'h4; //> 
    18'h12865: Data = 4'h4; //> 
    18'h12866: Data = 4'h4; //> 
    18'h12867: Data = 4'h4; //> 
    18'h12868: Data = 4'h6; //[ 
    18'h12869: Data = 4'h4; //> 
    18'h12870: Data = 4'h4; //> 
    18'h12871: Data = 4'h4; //> 
    18'h12872: Data = 4'h4; //> 
    18'h12873: Data = 4'h4; //> 
    18'h12874: Data = 4'h4; //> 
    18'h12875: Data = 4'h4; //> 
    18'h12876: Data = 4'h4; //> 
    18'h12877: Data = 4'h4; //> 
    18'h12878: Data = 4'h7; //] 
    18'h12879: Data = 4'h5; //< 
    18'h12880: Data = 4'h5; //< 
    18'h12881: Data = 4'h5; //< 
    18'h12882: Data = 4'h5; //< 
    18'h12883: Data = 4'h5; //< 
    18'h12884: Data = 4'h5; //< 
    18'h12885: Data = 4'h5; //< 
    18'h12886: Data = 4'h5; //< 
    18'h12887: Data = 4'h5; //< 
    18'h12888: Data = 4'h6; //[ 
    18'h12889: Data = 4'h4; //> 
    18'h12890: Data = 4'h6; //[ 
    18'h12891: Data = 4'h3; //- 
    18'h12892: Data = 4'h4; //> 
    18'h12893: Data = 4'h4; //> 
    18'h12894: Data = 4'h4; //> 
    18'h12895: Data = 4'h4; //> 
    18'h12896: Data = 4'h4; //> 
    18'h12897: Data = 4'h4; //> 
    18'h12898: Data = 4'h4; //> 
    18'h12899: Data = 4'h4; //> 
    18'h12900: Data = 4'h4; //> 
    18'h12901: Data = 4'h2; //+ 
    18'h12902: Data = 4'h5; //< 
    18'h12903: Data = 4'h5; //< 
    18'h12904: Data = 4'h5; //< 
    18'h12905: Data = 4'h5; //< 
    18'h12906: Data = 4'h5; //< 
    18'h12907: Data = 4'h5; //< 
    18'h12908: Data = 4'h5; //< 
    18'h12909: Data = 4'h5; //< 
    18'h12910: Data = 4'h5; //< 
    18'h12911: Data = 4'h7; //] 
    18'h12912: Data = 4'h5; //< 
    18'h12913: Data = 4'h5; //< 
    18'h12914: Data = 4'h5; //< 
    18'h12915: Data = 4'h5; //< 
    18'h12916: Data = 4'h5; //< 
    18'h12917: Data = 4'h5; //< 
    18'h12918: Data = 4'h5; //< 
    18'h12919: Data = 4'h5; //< 
    18'h12920: Data = 4'h5; //< 
    18'h12921: Data = 4'h5; //< 
    18'h12922: Data = 4'h7; //] 
    18'h12923: Data = 4'h4; //> 
    18'h12924: Data = 4'h6; //[ 
    18'h12925: Data = 4'h3; //- 
    18'h12926: Data = 4'h4; //> 
    18'h12927: Data = 4'h4; //> 
    18'h12928: Data = 4'h4; //> 
    18'h12929: Data = 4'h4; //> 
    18'h12930: Data = 4'h4; //> 
    18'h12931: Data = 4'h4; //> 
    18'h12932: Data = 4'h4; //> 
    18'h12933: Data = 4'h4; //> 
    18'h12934: Data = 4'h4; //> 
    18'h12935: Data = 4'h2; //+ 
    18'h12936: Data = 4'h5; //< 
    18'h12937: Data = 4'h5; //< 
    18'h12938: Data = 4'h5; //< 
    18'h12939: Data = 4'h5; //< 
    18'h12940: Data = 4'h5; //< 
    18'h12941: Data = 4'h5; //< 
    18'h12942: Data = 4'h5; //< 
    18'h12943: Data = 4'h5; //< 
    18'h12944: Data = 4'h5; //< 
    18'h12945: Data = 4'h7; //] 
    18'h12946: Data = 4'h5; //< 
    18'h12947: Data = 4'h2; //+ 
    18'h12948: Data = 4'h4; //> 
    18'h12949: Data = 4'h4; //> 
    18'h12950: Data = 4'h4; //> 
    18'h12951: Data = 4'h4; //> 
    18'h12952: Data = 4'h4; //> 
    18'h12953: Data = 4'h4; //> 
    18'h12954: Data = 4'h4; //> 
    18'h12955: Data = 4'h4; //> 
    18'h12956: Data = 4'h7; //] 
    18'h12957: Data = 4'h5; //< 
    18'h12958: Data = 4'h5; //< 
    18'h12959: Data = 4'h5; //< 
    18'h12960: Data = 4'h5; //< 
    18'h12961: Data = 4'h5; //< 
    18'h12962: Data = 4'h5; //< 
    18'h12963: Data = 4'h5; //< 
    18'h12964: Data = 4'h5; //< 
    18'h12965: Data = 4'h5; //< 
    18'h12966: Data = 4'h6; //[ 
    18'h12967: Data = 4'h4; //> 
    18'h12968: Data = 4'h6; //[ 
    18'h12969: Data = 4'h3; //- 
    18'h12970: Data = 4'h7; //] 
    18'h12971: Data = 4'h5; //< 
    18'h12972: Data = 4'h3; //- 
    18'h12973: Data = 4'h4; //> 
    18'h12974: Data = 4'h4; //> 
    18'h12975: Data = 4'h4; //> 
    18'h12976: Data = 4'h4; //> 
    18'h12977: Data = 4'h6; //[ 
    18'h12978: Data = 4'h3; //- 
    18'h12979: Data = 4'h5; //< 
    18'h12980: Data = 4'h5; //< 
    18'h12981: Data = 4'h5; //< 
    18'h12982: Data = 4'h5; //< 
    18'h12983: Data = 4'h2; //+ 
    18'h12984: Data = 4'h4; //> 
    18'h12985: Data = 4'h6; //[ 
    18'h12986: Data = 4'h5; //< 
    18'h12987: Data = 4'h3; //- 
    18'h12988: Data = 4'h4; //> 
    18'h12989: Data = 4'h3; //- 
    18'h12990: Data = 4'h5; //< 
    18'h12991: Data = 4'h5; //< 
    18'h12992: Data = 4'h5; //< 
    18'h12993: Data = 4'h5; //< 
    18'h12994: Data = 4'h5; //< 
    18'h12995: Data = 4'h5; //< 
    18'h12996: Data = 4'h2; //+ 
    18'h12997: Data = 4'h4; //> 
    18'h12998: Data = 4'h4; //> 
    18'h12999: Data = 4'h4; //> 
    18'h13000: Data = 4'h4; //> 
    18'h13001: Data = 4'h4; //> 
    18'h13002: Data = 4'h4; //> 
    18'h13003: Data = 4'h7; //] 
    18'h13004: Data = 4'h5; //< 
    18'h13005: Data = 4'h6; //[ 
    18'h13006: Data = 4'h3; //- 
    18'h13007: Data = 4'h4; //> 
    18'h13008: Data = 4'h2; //+ 
    18'h13009: Data = 4'h5; //< 
    18'h13010: Data = 4'h7; //] 
    18'h13011: Data = 4'h4; //> 
    18'h13012: Data = 4'h4; //> 
    18'h13013: Data = 4'h4; //> 
    18'h13014: Data = 4'h4; //> 
    18'h13015: Data = 4'h7; //] 
    18'h13016: Data = 4'h5; //< 
    18'h13017: Data = 4'h5; //< 
    18'h13018: Data = 4'h5; //< 
    18'h13019: Data = 4'h6; //[ 
    18'h13020: Data = 4'h3; //- 
    18'h13021: Data = 4'h4; //> 
    18'h13022: Data = 4'h4; //> 
    18'h13023: Data = 4'h4; //> 
    18'h13024: Data = 4'h2; //+ 
    18'h13025: Data = 4'h5; //< 
    18'h13026: Data = 4'h5; //< 
    18'h13027: Data = 4'h5; //< 
    18'h13028: Data = 4'h7; //] 
    18'h13029: Data = 4'h5; //< 
    18'h13030: Data = 4'h2; //+ 
    18'h13031: Data = 4'h5; //< 
    18'h13032: Data = 4'h5; //< 
    18'h13033: Data = 4'h5; //< 
    18'h13034: Data = 4'h5; //< 
    18'h13035: Data = 4'h5; //< 
    18'h13036: Data = 4'h5; //< 
    18'h13037: Data = 4'h5; //< 
    18'h13038: Data = 4'h5; //< 
    18'h13039: Data = 4'h5; //< 
    18'h13040: Data = 4'h7; //] 
    18'h13041: Data = 4'h4; //> 
    18'h13042: Data = 4'h4; //> 
    18'h13043: Data = 4'h4; //> 
    18'h13044: Data = 4'h4; //> 
    18'h13045: Data = 4'h4; //> 
    18'h13046: Data = 4'h4; //> 
    18'h13047: Data = 4'h4; //> 
    18'h13048: Data = 4'h4; //> 
    18'h13049: Data = 4'h4; //> 
    18'h13050: Data = 4'h6; //[ 
    18'h13051: Data = 4'h4; //> 
    18'h13052: Data = 4'h4; //> 
    18'h13053: Data = 4'h4; //> 
    18'h13054: Data = 4'h4; //> 
    18'h13055: Data = 4'h6; //[ 
    18'h13056: Data = 4'h3; //- 
    18'h13057: Data = 4'h5; //< 
    18'h13058: Data = 4'h5; //< 
    18'h13059: Data = 4'h5; //< 
    18'h13060: Data = 4'h5; //< 
    18'h13061: Data = 4'h5; //< 
    18'h13062: Data = 4'h5; //< 
    18'h13063: Data = 4'h5; //< 
    18'h13064: Data = 4'h5; //< 
    18'h13065: Data = 4'h5; //< 
    18'h13066: Data = 4'h5; //< 
    18'h13067: Data = 4'h5; //< 
    18'h13068: Data = 4'h5; //< 
    18'h13069: Data = 4'h5; //< 
    18'h13070: Data = 4'h5; //< 
    18'h13071: Data = 4'h5; //< 
    18'h13072: Data = 4'h5; //< 
    18'h13073: Data = 4'h5; //< 
    18'h13074: Data = 4'h5; //< 
    18'h13075: Data = 4'h5; //< 
    18'h13076: Data = 4'h5; //< 
    18'h13077: Data = 4'h5; //< 
    18'h13078: Data = 4'h5; //< 
    18'h13079: Data = 4'h5; //< 
    18'h13080: Data = 4'h5; //< 
    18'h13081: Data = 4'h5; //< 
    18'h13082: Data = 4'h5; //< 
    18'h13083: Data = 4'h5; //< 
    18'h13084: Data = 4'h5; //< 
    18'h13085: Data = 4'h5; //< 
    18'h13086: Data = 4'h5; //< 
    18'h13087: Data = 4'h5; //< 
    18'h13088: Data = 4'h5; //< 
    18'h13089: Data = 4'h5; //< 
    18'h13090: Data = 4'h5; //< 
    18'h13091: Data = 4'h5; //< 
    18'h13092: Data = 4'h5; //< 
    18'h13093: Data = 4'h2; //+ 
    18'h13094: Data = 4'h4; //> 
    18'h13095: Data = 4'h4; //> 
    18'h13096: Data = 4'h4; //> 
    18'h13097: Data = 4'h4; //> 
    18'h13098: Data = 4'h4; //> 
    18'h13099: Data = 4'h4; //> 
    18'h13100: Data = 4'h4; //> 
    18'h13101: Data = 4'h4; //> 
    18'h13102: Data = 4'h4; //> 
    18'h13103: Data = 4'h4; //> 
    18'h13104: Data = 4'h4; //> 
    18'h13105: Data = 4'h4; //> 
    18'h13106: Data = 4'h4; //> 
    18'h13107: Data = 4'h4; //> 
    18'h13108: Data = 4'h4; //> 
    18'h13109: Data = 4'h4; //> 
    18'h13110: Data = 4'h4; //> 
    18'h13111: Data = 4'h4; //> 
    18'h13112: Data = 4'h4; //> 
    18'h13113: Data = 4'h4; //> 
    18'h13114: Data = 4'h4; //> 
    18'h13115: Data = 4'h4; //> 
    18'h13116: Data = 4'h4; //> 
    18'h13117: Data = 4'h4; //> 
    18'h13118: Data = 4'h4; //> 
    18'h13119: Data = 4'h4; //> 
    18'h13120: Data = 4'h4; //> 
    18'h13121: Data = 4'h4; //> 
    18'h13122: Data = 4'h4; //> 
    18'h13123: Data = 4'h4; //> 
    18'h13124: Data = 4'h4; //> 
    18'h13125: Data = 4'h4; //> 
    18'h13126: Data = 4'h4; //> 
    18'h13127: Data = 4'h4; //> 
    18'h13128: Data = 4'h4; //> 
    18'h13129: Data = 4'h4; //> 
    18'h13130: Data = 4'h7; //] 
    18'h13131: Data = 4'h4; //> 
    18'h13132: Data = 4'h4; //> 
    18'h13133: Data = 4'h4; //> 
    18'h13134: Data = 4'h4; //> 
    18'h13135: Data = 4'h4; //> 
    18'h13136: Data = 4'h7; //] 
    18'h13137: Data = 4'h5; //< 
    18'h13138: Data = 4'h5; //< 
    18'h13139: Data = 4'h5; //< 
    18'h13140: Data = 4'h5; //< 
    18'h13141: Data = 4'h5; //< 
    18'h13142: Data = 4'h5; //< 
    18'h13143: Data = 4'h5; //< 
    18'h13144: Data = 4'h5; //< 
    18'h13145: Data = 4'h5; //< 
    18'h13146: Data = 4'h6; //[ 
    18'h13147: Data = 4'h5; //< 
    18'h13148: Data = 4'h5; //< 
    18'h13149: Data = 4'h5; //< 
    18'h13150: Data = 4'h5; //< 
    18'h13151: Data = 4'h5; //< 
    18'h13152: Data = 4'h5; //< 
    18'h13153: Data = 4'h5; //< 
    18'h13154: Data = 4'h5; //< 
    18'h13155: Data = 4'h5; //< 
    18'h13156: Data = 4'h7; //] 
    18'h13157: Data = 4'h4; //> 
    18'h13158: Data = 4'h4; //> 
    18'h13159: Data = 4'h4; //> 
    18'h13160: Data = 4'h4; //> 
    18'h13161: Data = 4'h4; //> 
    18'h13162: Data = 4'h4; //> 
    18'h13163: Data = 4'h4; //> 
    18'h13164: Data = 4'h4; //> 
    18'h13165: Data = 4'h4; //> 
    18'h13166: Data = 4'h6; //[ 
    18'h13167: Data = 4'h4; //> 
    18'h13168: Data = 4'h4; //> 
    18'h13169: Data = 4'h4; //> 
    18'h13170: Data = 4'h6; //[ 
    18'h13171: Data = 4'h3; //- 
    18'h13172: Data = 4'h5; //< 
    18'h13173: Data = 4'h5; //< 
    18'h13174: Data = 4'h5; //< 
    18'h13175: Data = 4'h5; //< 
    18'h13176: Data = 4'h5; //< 
    18'h13177: Data = 4'h5; //< 
    18'h13178: Data = 4'h5; //< 
    18'h13179: Data = 4'h5; //< 
    18'h13180: Data = 4'h5; //< 
    18'h13181: Data = 4'h5; //< 
    18'h13182: Data = 4'h5; //< 
    18'h13183: Data = 4'h5; //< 
    18'h13184: Data = 4'h5; //< 
    18'h13185: Data = 4'h5; //< 
    18'h13186: Data = 4'h5; //< 
    18'h13187: Data = 4'h5; //< 
    18'h13188: Data = 4'h5; //< 
    18'h13189: Data = 4'h5; //< 
    18'h13190: Data = 4'h5; //< 
    18'h13191: Data = 4'h5; //< 
    18'h13192: Data = 4'h5; //< 
    18'h13193: Data = 4'h5; //< 
    18'h13194: Data = 4'h5; //< 
    18'h13195: Data = 4'h5; //< 
    18'h13196: Data = 4'h5; //< 
    18'h13197: Data = 4'h5; //< 
    18'h13198: Data = 4'h5; //< 
    18'h13199: Data = 4'h5; //< 
    18'h13200: Data = 4'h5; //< 
    18'h13201: Data = 4'h5; //< 
    18'h13202: Data = 4'h5; //< 
    18'h13203: Data = 4'h5; //< 
    18'h13204: Data = 4'h5; //< 
    18'h13205: Data = 4'h5; //< 
    18'h13206: Data = 4'h5; //< 
    18'h13207: Data = 4'h5; //< 
    18'h13208: Data = 4'h2; //+ 
    18'h13209: Data = 4'h4; //> 
    18'h13210: Data = 4'h4; //> 
    18'h13211: Data = 4'h4; //> 
    18'h13212: Data = 4'h4; //> 
    18'h13213: Data = 4'h4; //> 
    18'h13214: Data = 4'h4; //> 
    18'h13215: Data = 4'h4; //> 
    18'h13216: Data = 4'h4; //> 
    18'h13217: Data = 4'h4; //> 
    18'h13218: Data = 4'h4; //> 
    18'h13219: Data = 4'h4; //> 
    18'h13220: Data = 4'h4; //> 
    18'h13221: Data = 4'h4; //> 
    18'h13222: Data = 4'h4; //> 
    18'h13223: Data = 4'h4; //> 
    18'h13224: Data = 4'h4; //> 
    18'h13225: Data = 4'h4; //> 
    18'h13226: Data = 4'h4; //> 
    18'h13227: Data = 4'h4; //> 
    18'h13228: Data = 4'h4; //> 
    18'h13229: Data = 4'h4; //> 
    18'h13230: Data = 4'h4; //> 
    18'h13231: Data = 4'h4; //> 
    18'h13232: Data = 4'h4; //> 
    18'h13233: Data = 4'h4; //> 
    18'h13234: Data = 4'h4; //> 
    18'h13235: Data = 4'h4; //> 
    18'h13236: Data = 4'h4; //> 
    18'h13237: Data = 4'h4; //> 
    18'h13238: Data = 4'h4; //> 
    18'h13239: Data = 4'h4; //> 
    18'h13240: Data = 4'h4; //> 
    18'h13241: Data = 4'h4; //> 
    18'h13242: Data = 4'h4; //> 
    18'h13243: Data = 4'h4; //> 
    18'h13244: Data = 4'h4; //> 
    18'h13245: Data = 4'h7; //] 
    18'h13246: Data = 4'h4; //> 
    18'h13247: Data = 4'h4; //> 
    18'h13248: Data = 4'h4; //> 
    18'h13249: Data = 4'h4; //> 
    18'h13250: Data = 4'h4; //> 
    18'h13251: Data = 4'h4; //> 
    18'h13252: Data = 4'h7; //] 
    18'h13253: Data = 4'h5; //< 
    18'h13254: Data = 4'h5; //< 
    18'h13255: Data = 4'h5; //< 
    18'h13256: Data = 4'h5; //< 
    18'h13257: Data = 4'h5; //< 
    18'h13258: Data = 4'h5; //< 
    18'h13259: Data = 4'h5; //< 
    18'h13260: Data = 4'h5; //< 
    18'h13261: Data = 4'h5; //< 
    18'h13262: Data = 4'h6; //[ 
    18'h13263: Data = 4'h5; //< 
    18'h13264: Data = 4'h5; //< 
    18'h13265: Data = 4'h5; //< 
    18'h13266: Data = 4'h5; //< 
    18'h13267: Data = 4'h5; //< 
    18'h13268: Data = 4'h5; //< 
    18'h13269: Data = 4'h5; //< 
    18'h13270: Data = 4'h5; //< 
    18'h13271: Data = 4'h5; //< 
    18'h13272: Data = 4'h7; //] 
    18'h13273: Data = 4'h4; //> 
    18'h13274: Data = 4'h4; //> 
    18'h13275: Data = 4'h4; //> 
    18'h13276: Data = 4'h4; //> 
    18'h13277: Data = 4'h4; //> 
    18'h13278: Data = 4'h4; //> 
    18'h13279: Data = 4'h4; //> 
    18'h13280: Data = 4'h4; //> 
    18'h13281: Data = 4'h4; //> 
    18'h13282: Data = 4'h2; //+ 
    18'h13283: Data = 4'h2; //+ 
    18'h13284: Data = 4'h2; //+ 
    18'h13285: Data = 4'h2; //+ 
    18'h13286: Data = 4'h2; //+ 
    18'h13287: Data = 4'h2; //+ 
    18'h13288: Data = 4'h2; //+ 
    18'h13289: Data = 4'h2; //+ 
    18'h13290: Data = 4'h2; //+ 
    18'h13291: Data = 4'h2; //+ 
    18'h13292: Data = 4'h2; //+ 
    18'h13293: Data = 4'h2; //+ 
    18'h13294: Data = 4'h2; //+ 
    18'h13295: Data = 4'h2; //+ 
    18'h13296: Data = 4'h2; //+ 
    18'h13297: Data = 4'h6; //[ 
    18'h13298: Data = 4'h6; //[ 
    18'h13299: Data = 4'h4; //> 
    18'h13300: Data = 4'h4; //> 
    18'h13301: Data = 4'h4; //> 
    18'h13302: Data = 4'h4; //> 
    18'h13303: Data = 4'h4; //> 
    18'h13304: Data = 4'h4; //> 
    18'h13305: Data = 4'h4; //> 
    18'h13306: Data = 4'h4; //> 
    18'h13307: Data = 4'h4; //> 
    18'h13308: Data = 4'h7; //] 
    18'h13309: Data = 4'h5; //< 
    18'h13310: Data = 4'h5; //< 
    18'h13311: Data = 4'h5; //< 
    18'h13312: Data = 4'h5; //< 
    18'h13313: Data = 4'h5; //< 
    18'h13314: Data = 4'h5; //< 
    18'h13315: Data = 4'h5; //< 
    18'h13316: Data = 4'h5; //< 
    18'h13317: Data = 4'h5; //< 
    18'h13318: Data = 4'h3; //- 
    18'h13319: Data = 4'h5; //< 
    18'h13320: Data = 4'h5; //< 
    18'h13321: Data = 4'h5; //< 
    18'h13322: Data = 4'h5; //< 
    18'h13323: Data = 4'h5; //< 
    18'h13324: Data = 4'h5; //< 
    18'h13325: Data = 4'h5; //< 
    18'h13326: Data = 4'h5; //< 
    18'h13327: Data = 4'h5; //< 
    18'h13328: Data = 4'h6; //[ 
    18'h13329: Data = 4'h5; //< 
    18'h13330: Data = 4'h5; //< 
    18'h13331: Data = 4'h5; //< 
    18'h13332: Data = 4'h5; //< 
    18'h13333: Data = 4'h5; //< 
    18'h13334: Data = 4'h5; //< 
    18'h13335: Data = 4'h5; //< 
    18'h13336: Data = 4'h5; //< 
    18'h13337: Data = 4'h5; //< 
    18'h13338: Data = 4'h7; //] 
    18'h13339: Data = 4'h4; //> 
    18'h13340: Data = 4'h4; //> 
    18'h13341: Data = 4'h4; //> 
    18'h13342: Data = 4'h4; //> 
    18'h13343: Data = 4'h4; //> 
    18'h13344: Data = 4'h4; //> 
    18'h13345: Data = 4'h4; //> 
    18'h13346: Data = 4'h4; //> 
    18'h13347: Data = 4'h4; //> 
    18'h13348: Data = 4'h3; //- 
    18'h13349: Data = 4'h7; //] 
    18'h13350: Data = 4'h2; //+ 
    18'h13351: Data = 4'h6; //[ 
    18'h13352: Data = 4'h4; //> 
    18'h13353: Data = 4'h4; //> 
    18'h13354: Data = 4'h4; //> 
    18'h13355: Data = 4'h4; //> 
    18'h13356: Data = 4'h4; //> 
    18'h13357: Data = 4'h4; //> 
    18'h13358: Data = 4'h4; //> 
    18'h13359: Data = 4'h4; //> 
    18'h13360: Data = 4'h6; //[ 
    18'h13361: Data = 4'h3; //- 
    18'h13362: Data = 4'h5; //< 
    18'h13363: Data = 4'h5; //< 
    18'h13364: Data = 4'h5; //< 
    18'h13365: Data = 4'h5; //< 
    18'h13366: Data = 4'h5; //< 
    18'h13367: Data = 4'h5; //< 
    18'h13368: Data = 4'h5; //< 
    18'h13369: Data = 4'h2; //+ 
    18'h13370: Data = 4'h4; //> 
    18'h13371: Data = 4'h4; //> 
    18'h13372: Data = 4'h4; //> 
    18'h13373: Data = 4'h4; //> 
    18'h13374: Data = 4'h4; //> 
    18'h13375: Data = 4'h4; //> 
    18'h13376: Data = 4'h4; //> 
    18'h13377: Data = 4'h7; //] 
    18'h13378: Data = 4'h5; //< 
    18'h13379: Data = 4'h5; //< 
    18'h13380: Data = 4'h5; //< 
    18'h13381: Data = 4'h5; //< 
    18'h13382: Data = 4'h5; //< 
    18'h13383: Data = 4'h5; //< 
    18'h13384: Data = 4'h5; //< 
    18'h13385: Data = 4'h6; //[ 
    18'h13386: Data = 4'h3; //- 
    18'h13387: Data = 4'h4; //> 
    18'h13388: Data = 4'h4; //> 
    18'h13389: Data = 4'h4; //> 
    18'h13390: Data = 4'h4; //> 
    18'h13391: Data = 4'h4; //> 
    18'h13392: Data = 4'h4; //> 
    18'h13393: Data = 4'h4; //> 
    18'h13394: Data = 4'h2; //+ 
    18'h13395: Data = 4'h5; //< 
    18'h13396: Data = 4'h5; //< 
    18'h13397: Data = 4'h5; //< 
    18'h13398: Data = 4'h5; //< 
    18'h13399: Data = 4'h5; //< 
    18'h13400: Data = 4'h5; //< 
    18'h13401: Data = 4'h2; //+ 
    18'h13402: Data = 4'h5; //< 
    18'h13403: Data = 4'h7; //] 
    18'h13404: Data = 4'h4; //> 
    18'h13405: Data = 4'h4; //> 
    18'h13406: Data = 4'h4; //> 
    18'h13407: Data = 4'h4; //> 
    18'h13408: Data = 4'h4; //> 
    18'h13409: Data = 4'h4; //> 
    18'h13410: Data = 4'h4; //> 
    18'h13411: Data = 4'h4; //> 
    18'h13412: Data = 4'h7; //] 
    18'h13413: Data = 4'h5; //< 
    18'h13414: Data = 4'h5; //< 
    18'h13415: Data = 4'h5; //< 
    18'h13416: Data = 4'h5; //< 
    18'h13417: Data = 4'h5; //< 
    18'h13418: Data = 4'h5; //< 
    18'h13419: Data = 4'h5; //< 
    18'h13420: Data = 4'h5; //< 
    18'h13421: Data = 4'h5; //< 
    18'h13422: Data = 4'h6; //[ 
    18'h13423: Data = 4'h5; //< 
    18'h13424: Data = 4'h5; //< 
    18'h13425: Data = 4'h5; //< 
    18'h13426: Data = 4'h5; //< 
    18'h13427: Data = 4'h5; //< 
    18'h13428: Data = 4'h5; //< 
    18'h13429: Data = 4'h5; //< 
    18'h13430: Data = 4'h5; //< 
    18'h13431: Data = 4'h5; //< 
    18'h13432: Data = 4'h7; //] 
    18'h13433: Data = 4'h4; //> 
    18'h13434: Data = 4'h4; //> 
    18'h13435: Data = 4'h4; //> 
    18'h13436: Data = 4'h4; //> 
    18'h13437: Data = 4'h4; //> 
    18'h13438: Data = 4'h4; //> 
    18'h13439: Data = 4'h4; //> 
    18'h13440: Data = 4'h4; //> 
    18'h13441: Data = 4'h4; //> 
    18'h13442: Data = 4'h6; //[ 
    18'h13443: Data = 4'h4; //> 
    18'h13444: Data = 4'h4; //> 
    18'h13445: Data = 4'h4; //> 
    18'h13446: Data = 4'h4; //> 
    18'h13447: Data = 4'h4; //> 
    18'h13448: Data = 4'h4; //> 
    18'h13449: Data = 4'h6; //[ 
    18'h13450: Data = 4'h3; //- 
    18'h13451: Data = 4'h7; //] 
    18'h13452: Data = 4'h4; //> 
    18'h13453: Data = 4'h4; //> 
    18'h13454: Data = 4'h4; //> 
    18'h13455: Data = 4'h7; //] 
    18'h13456: Data = 4'h5; //< 
    18'h13457: Data = 4'h5; //< 
    18'h13458: Data = 4'h5; //< 
    18'h13459: Data = 4'h5; //< 
    18'h13460: Data = 4'h5; //< 
    18'h13461: Data = 4'h5; //< 
    18'h13462: Data = 4'h5; //< 
    18'h13463: Data = 4'h5; //< 
    18'h13464: Data = 4'h5; //< 
    18'h13465: Data = 4'h6; //[ 
    18'h13466: Data = 4'h5; //< 
    18'h13467: Data = 4'h5; //< 
    18'h13468: Data = 4'h5; //< 
    18'h13469: Data = 4'h5; //< 
    18'h13470: Data = 4'h5; //< 
    18'h13471: Data = 4'h5; //< 
    18'h13472: Data = 4'h5; //< 
    18'h13473: Data = 4'h5; //< 
    18'h13474: Data = 4'h5; //< 
    18'h13475: Data = 4'h7; //] 
    18'h13476: Data = 4'h4; //> 
    18'h13477: Data = 4'h4; //> 
    18'h13478: Data = 4'h4; //> 
    18'h13479: Data = 4'h4; //> 
    18'h13480: Data = 4'h2; //+ 
    18'h13481: Data = 4'h4; //> 
    18'h13482: Data = 4'h6; //[ 
    18'h13483: Data = 4'h3; //- 
    18'h13484: Data = 4'h5; //< 
    18'h13485: Data = 4'h3; //- 
    18'h13486: Data = 4'h5; //< 
    18'h13487: Data = 4'h5; //< 
    18'h13488: Data = 4'h5; //< 
    18'h13489: Data = 4'h5; //< 
    18'h13490: Data = 4'h2; //+ 
    18'h13491: Data = 4'h4; //> 
    18'h13492: Data = 4'h4; //> 
    18'h13493: Data = 4'h4; //> 
    18'h13494: Data = 4'h4; //> 
    18'h13495: Data = 4'h4; //> 
    18'h13496: Data = 4'h7; //] 
    18'h13497: Data = 4'h4; //> 
    18'h13498: Data = 4'h6; //[ 
    18'h13499: Data = 4'h3; //- 
    18'h13500: Data = 4'h5; //< 
    18'h13501: Data = 4'h5; //< 
    18'h13502: Data = 4'h5; //< 
    18'h13503: Data = 4'h5; //< 
    18'h13504: Data = 4'h5; //< 
    18'h13505: Data = 4'h5; //< 
    18'h13506: Data = 4'h6; //[ 
    18'h13507: Data = 4'h3; //- 
    18'h13508: Data = 4'h4; //> 
    18'h13509: Data = 4'h4; //> 
    18'h13510: Data = 4'h4; //> 
    18'h13511: Data = 4'h4; //> 
    18'h13512: Data = 4'h4; //> 
    18'h13513: Data = 4'h2; //+ 
    18'h13514: Data = 4'h5; //< 
    18'h13515: Data = 4'h2; //+ 
    18'h13516: Data = 4'h2; //+ 
    18'h13517: Data = 4'h5; //< 
    18'h13518: Data = 4'h5; //< 
    18'h13519: Data = 4'h5; //< 
    18'h13520: Data = 4'h5; //< 
    18'h13521: Data = 4'h7; //] 
    18'h13522: Data = 4'h4; //> 
    18'h13523: Data = 4'h4; //> 
    18'h13524: Data = 4'h4; //> 
    18'h13525: Data = 4'h4; //> 
    18'h13526: Data = 4'h4; //> 
    18'h13527: Data = 4'h6; //[ 
    18'h13528: Data = 4'h3; //- 
    18'h13529: Data = 4'h5; //< 
    18'h13530: Data = 4'h5; //< 
    18'h13531: Data = 4'h5; //< 
    18'h13532: Data = 4'h5; //< 
    18'h13533: Data = 4'h5; //< 
    18'h13534: Data = 4'h2; //+ 
    18'h13535: Data = 4'h4; //> 
    18'h13536: Data = 4'h4; //> 
    18'h13537: Data = 4'h4; //> 
    18'h13538: Data = 4'h4; //> 
    18'h13539: Data = 4'h4; //> 
    18'h13540: Data = 4'h7; //] 
    18'h13541: Data = 4'h5; //< 
    18'h13542: Data = 4'h3; //- 
    18'h13543: Data = 4'h4; //> 
    18'h13544: Data = 4'h2; //+ 
    18'h13545: Data = 4'h4; //> 
    18'h13546: Data = 4'h7; //] 
    18'h13547: Data = 4'h5; //< 
    18'h13548: Data = 4'h6; //[ 
    18'h13549: Data = 4'h3; //- 
    18'h13550: Data = 4'h4; //> 
    18'h13551: Data = 4'h2; //+ 
    18'h13552: Data = 4'h5; //< 
    18'h13553: Data = 4'h7; //] 
    18'h13554: Data = 4'h5; //< 
    18'h13555: Data = 4'h5; //< 
    18'h13556: Data = 4'h5; //< 
    18'h13557: Data = 4'h5; //< 
    18'h13558: Data = 4'h5; //< 
    18'h13559: Data = 4'h6; //[ 
    18'h13560: Data = 4'h3; //- 
    18'h13561: Data = 4'h4; //> 
    18'h13562: Data = 4'h4; //> 
    18'h13563: Data = 4'h4; //> 
    18'h13564: Data = 4'h4; //> 
    18'h13565: Data = 4'h4; //> 
    18'h13566: Data = 4'h2; //+ 
    18'h13567: Data = 4'h5; //< 
    18'h13568: Data = 4'h5; //< 
    18'h13569: Data = 4'h5; //< 
    18'h13570: Data = 4'h5; //< 
    18'h13571: Data = 4'h5; //< 
    18'h13572: Data = 4'h7; //] 
    18'h13573: Data = 4'h4; //> 
    18'h13574: Data = 4'h4; //> 
    18'h13575: Data = 4'h4; //> 
    18'h13576: Data = 4'h4; //> 
    18'h13577: Data = 4'h4; //> 
    18'h13578: Data = 4'h4; //> 
    18'h13579: Data = 4'ha; //0 
    18'h13580: Data = 4'h5; //< 
    18'h13581: Data = 4'h5; //< 
    18'h13582: Data = 4'h5; //< 
    18'h13583: Data = 4'h5; //< 
    18'h13584: Data = 4'h5; //< 
    18'h13585: Data = 4'h5; //< 
    18'h13586: Data = 4'h2; //+ 
    18'h13587: Data = 4'h4; //> 
    18'h13588: Data = 4'h4; //> 
    18'h13589: Data = 4'h4; //> 
    18'h13590: Data = 4'h4; //> 
    18'h13591: Data = 4'h6; //[ 
    18'h13592: Data = 4'h3; //- 
    18'h13593: Data = 4'h5; //< 
    18'h13594: Data = 4'h5; //< 
    18'h13595: Data = 4'h5; //< 
    18'h13596: Data = 4'h5; //< 
    18'h13597: Data = 4'h3; //- 
    18'h13598: Data = 4'h4; //> 
    18'h13599: Data = 4'h4; //> 
    18'h13600: Data = 4'h4; //> 
    18'h13601: Data = 4'h4; //> 
    18'h13602: Data = 4'h7; //] 
    18'h13603: Data = 4'h2; //+ 
    18'h13604: Data = 4'h5; //< 
    18'h13605: Data = 4'h5; //< 
    18'h13606: Data = 4'h5; //< 
    18'h13607: Data = 4'h5; //< 
    18'h13608: Data = 4'h6; //[ 
    18'h13609: Data = 4'h3; //- 
    18'h13610: Data = 4'h4; //> 
    18'h13611: Data = 4'h4; //> 
    18'h13612: Data = 4'h4; //> 
    18'h13613: Data = 4'h4; //> 
    18'h13614: Data = 4'h3; //- 
    18'h13615: Data = 4'h4; //> 
    18'h13616: Data = 4'h4; //> 
    18'h13617: Data = 4'h4; //> 
    18'h13618: Data = 4'h4; //> 
    18'h13619: Data = 4'h4; //> 
    18'h13620: Data = 4'h6; //[ 
    18'h13621: Data = 4'h4; //> 
    18'h13622: Data = 4'h4; //> 
    18'h13623: Data = 4'h6; //[ 
    18'h13624: Data = 4'h3; //- 
    18'h13625: Data = 4'h5; //< 
    18'h13626: Data = 4'h5; //< 
    18'h13627: Data = 4'h3; //- 
    18'h13628: Data = 4'h4; //> 
    18'h13629: Data = 4'h4; //> 
    18'h13630: Data = 4'h7; //] 
    18'h13631: Data = 4'h2; //+ 
    18'h13632: Data = 4'h5; //< 
    18'h13633: Data = 4'h5; //< 
    18'h13634: Data = 4'h6; //[ 
    18'h13635: Data = 4'h3; //- 
    18'h13636: Data = 4'h4; //> 
    18'h13637: Data = 4'h4; //> 
    18'h13638: Data = 4'h3; //- 
    18'h13639: Data = 4'h4; //> 
    18'h13640: Data = 4'h6; //[ 
    18'h13641: Data = 4'h3; //- 
    18'h13642: Data = 4'h5; //< 
    18'h13643: Data = 4'h5; //< 
    18'h13644: Data = 4'h5; //< 
    18'h13645: Data = 4'h2; //+ 
    18'h13646: Data = 4'h4; //> 
    18'h13647: Data = 4'h4; //> 
    18'h13648: Data = 4'h4; //> 
    18'h13649: Data = 4'h7; //] 
    18'h13650: Data = 4'h5; //< 
    18'h13651: Data = 4'h5; //< 
    18'h13652: Data = 4'h5; //< 
    18'h13653: Data = 4'h6; //[ 
    18'h13654: Data = 4'h3; //- 
    18'h13655: Data = 4'h4; //> 
    18'h13656: Data = 4'h4; //> 
    18'h13657: Data = 4'h4; //> 
    18'h13658: Data = 4'h2; //+ 
    18'h13659: Data = 4'h5; //< 
    18'h13660: Data = 4'h5; //< 
    18'h13661: Data = 4'h5; //< 
    18'h13662: Data = 4'h5; //< 
    18'h13663: Data = 4'h5; //< 
    18'h13664: Data = 4'h5; //< 
    18'h13665: Data = 4'h5; //< 
    18'h13666: Data = 4'h5; //< 
    18'h13667: Data = 4'h5; //< 
    18'h13668: Data = 4'h5; //< 
    18'h13669: Data = 4'h5; //< 
    18'h13670: Data = 4'h5; //< 
    18'h13671: Data = 4'h6; //[ 
    18'h13672: Data = 4'h5; //< 
    18'h13673: Data = 4'h5; //< 
    18'h13674: Data = 4'h5; //< 
    18'h13675: Data = 4'h5; //< 
    18'h13676: Data = 4'h5; //< 
    18'h13677: Data = 4'h5; //< 
    18'h13678: Data = 4'h5; //< 
    18'h13679: Data = 4'h5; //< 
    18'h13680: Data = 4'h5; //< 
    18'h13681: Data = 4'h7; //] 
    18'h13682: Data = 4'h4; //> 
    18'h13683: Data = 4'h4; //> 
    18'h13684: Data = 4'h4; //> 
    18'h13685: Data = 4'ha; //0 
    18'h13686: Data = 4'h2; //+ 
    18'h13687: Data = 4'h4; //> 
    18'h13688: Data = 4'h4; //> 
    18'h13689: Data = 4'h4; //> 
    18'h13690: Data = 4'h4; //> 
    18'h13691: Data = 4'h4; //> 
    18'h13692: Data = 4'h4; //> 
    18'h13693: Data = 4'h6; //[ 
    18'h13694: Data = 4'h4; //> 
    18'h13695: Data = 4'h4; //> 
    18'h13696: Data = 4'h4; //> 
    18'h13697: Data = 4'h4; //> 
    18'h13698: Data = 4'h4; //> 
    18'h13699: Data = 4'h4; //> 
    18'h13700: Data = 4'h4; //> 
    18'h13701: Data = 4'h4; //> 
    18'h13702: Data = 4'h4; //> 
    18'h13703: Data = 4'h7; //] 
    18'h13704: Data = 4'h4; //> 
    18'h13705: Data = 4'h2; //+ 
    18'h13706: Data = 4'h5; //< 
    18'h13707: Data = 4'h7; //] 
    18'h13708: Data = 4'h7; //] 
    18'h13709: Data = 4'h2; //+ 
    18'h13710: Data = 4'h4; //> 
    18'h13711: Data = 4'h4; //> 
    18'h13712: Data = 4'h4; //> 
    18'h13713: Data = 4'h6; //[ 
    18'h13714: Data = 4'h3; //- 
    18'h13715: Data = 4'h5; //< 
    18'h13716: Data = 4'h5; //< 
    18'h13717: Data = 4'h5; //< 
    18'h13718: Data = 4'h3; //- 
    18'h13719: Data = 4'h4; //> 
    18'h13720: Data = 4'h4; //> 
    18'h13721: Data = 4'h4; //> 
    18'h13722: Data = 4'h7; //] 
    18'h13723: Data = 4'h2; //+ 
    18'h13724: Data = 4'h5; //< 
    18'h13725: Data = 4'h5; //< 
    18'h13726: Data = 4'h5; //< 
    18'h13727: Data = 4'h6; //[ 
    18'h13728: Data = 4'h3; //- 
    18'h13729: Data = 4'h4; //> 
    18'h13730: Data = 4'h4; //> 
    18'h13731: Data = 4'h4; //> 
    18'h13732: Data = 4'h3; //- 
    18'h13733: Data = 4'h5; //< 
    18'h13734: Data = 4'h6; //[ 
    18'h13735: Data = 4'h3; //- 
    18'h13736: Data = 4'h5; //< 
    18'h13737: Data = 4'h5; //< 
    18'h13738: Data = 4'h2; //+ 
    18'h13739: Data = 4'h4; //> 
    18'h13740: Data = 4'h4; //> 
    18'h13741: Data = 4'h7; //] 
    18'h13742: Data = 4'h5; //< 
    18'h13743: Data = 4'h5; //< 
    18'h13744: Data = 4'h6; //[ 
    18'h13745: Data = 4'h3; //- 
    18'h13746: Data = 4'h4; //> 
    18'h13747: Data = 4'h4; //> 
    18'h13748: Data = 4'h2; //+ 
    18'h13749: Data = 4'h5; //< 
    18'h13750: Data = 4'h5; //< 
    18'h13751: Data = 4'h5; //< 
    18'h13752: Data = 4'h5; //< 
    18'h13753: Data = 4'h5; //< 
    18'h13754: Data = 4'h5; //< 
    18'h13755: Data = 4'h5; //< 
    18'h13756: Data = 4'h5; //< 
    18'h13757: Data = 4'h5; //< 
    18'h13758: Data = 4'h5; //< 
    18'h13759: Data = 4'h5; //< 
    18'h13760: Data = 4'h6; //[ 
    18'h13761: Data = 4'h5; //< 
    18'h13762: Data = 4'h5; //< 
    18'h13763: Data = 4'h5; //< 
    18'h13764: Data = 4'h5; //< 
    18'h13765: Data = 4'h5; //< 
    18'h13766: Data = 4'h5; //< 
    18'h13767: Data = 4'h5; //< 
    18'h13768: Data = 4'h5; //< 
    18'h13769: Data = 4'h5; //< 
    18'h13770: Data = 4'h7; //] 
    18'h13771: Data = 4'h4; //> 
    18'h13772: Data = 4'h4; //> 
    18'h13773: Data = 4'h4; //> 
    18'h13774: Data = 4'h4; //> 
    18'h13775: Data = 4'ha; //0 
    18'h13776: Data = 4'h2; //+ 
    18'h13777: Data = 4'h4; //> 
    18'h13778: Data = 4'h4; //> 
    18'h13779: Data = 4'h4; //> 
    18'h13780: Data = 4'h4; //> 
    18'h13781: Data = 4'h4; //> 
    18'h13782: Data = 4'h6; //[ 
    18'h13783: Data = 4'h4; //> 
    18'h13784: Data = 4'h4; //> 
    18'h13785: Data = 4'h4; //> 
    18'h13786: Data = 4'h4; //> 
    18'h13787: Data = 4'h4; //> 
    18'h13788: Data = 4'h4; //> 
    18'h13789: Data = 4'h4; //> 
    18'h13790: Data = 4'h4; //> 
    18'h13791: Data = 4'h4; //> 
    18'h13792: Data = 4'h7; //] 
    18'h13793: Data = 4'h4; //> 
    18'h13794: Data = 4'ha; //0 
    18'h13795: Data = 4'h2; //+ 
    18'h13796: Data = 4'h5; //< 
    18'h13797: Data = 4'h7; //] 
    18'h13798: Data = 4'h7; //] 
    18'h13799: Data = 4'h2; //+ 
    18'h13800: Data = 4'h4; //> 
    18'h13801: Data = 4'h6; //[ 
    18'h13802: Data = 4'h3; //- 
    18'h13803: Data = 4'h5; //< 
    18'h13804: Data = 4'h6; //[ 
    18'h13805: Data = 4'h4; //> 
    18'h13806: Data = 4'h4; //> 
    18'h13807: Data = 4'h4; //> 
    18'h13808: Data = 4'h4; //> 
    18'h13809: Data = 4'h4; //> 
    18'h13810: Data = 4'h4; //> 
    18'h13811: Data = 4'h4; //> 
    18'h13812: Data = 4'h4; //> 
    18'h13813: Data = 4'h4; //> 
    18'h13814: Data = 4'h7; //] 
    18'h13815: Data = 4'h5; //< 
    18'h13816: Data = 4'h5; //< 
    18'h13817: Data = 4'h5; //< 
    18'h13818: Data = 4'h5; //< 
    18'h13819: Data = 4'h5; //< 
    18'h13820: Data = 4'h5; //< 
    18'h13821: Data = 4'h5; //< 
    18'h13822: Data = 4'h5; //< 
    18'h13823: Data = 4'h7; //] 
    18'h13824: Data = 4'h4; //> 
    18'h13825: Data = 4'h4; //> 
    18'h13826: Data = 4'h4; //> 
    18'h13827: Data = 4'h4; //> 
    18'h13828: Data = 4'h4; //> 
    18'h13829: Data = 4'h4; //> 
    18'h13830: Data = 4'h4; //> 
    18'h13831: Data = 4'h4; //> 
    18'h13832: Data = 4'h7; //] 
    18'h13833: Data = 4'h5; //< 
    18'h13834: Data = 4'h5; //< 
    18'h13835: Data = 4'h5; //< 
    18'h13836: Data = 4'h5; //< 
    18'h13837: Data = 4'h5; //< 
    18'h13838: Data = 4'h5; //< 
    18'h13839: Data = 4'h5; //< 
    18'h13840: Data = 4'h5; //< 
    18'h13841: Data = 4'h5; //< 
    18'h13842: Data = 4'h6; //[ 
    18'h13843: Data = 4'h5; //< 
    18'h13844: Data = 4'h5; //< 
    18'h13845: Data = 4'h5; //< 
    18'h13846: Data = 4'h5; //< 
    18'h13847: Data = 4'h5; //< 
    18'h13848: Data = 4'h5; //< 
    18'h13849: Data = 4'h5; //< 
    18'h13850: Data = 4'h5; //< 
    18'h13851: Data = 4'h5; //< 
    18'h13852: Data = 4'h7; //] 
    18'h13853: Data = 4'h4; //> 
    18'h13854: Data = 4'h4; //> 
    18'h13855: Data = 4'h4; //> 
    18'h13856: Data = 4'h4; //> 
    18'h13857: Data = 4'h6; //[ 
    18'h13858: Data = 4'h3; //- 
    18'h13859: Data = 4'h5; //< 
    18'h13860: Data = 4'h5; //< 
    18'h13861: Data = 4'h5; //< 
    18'h13862: Data = 4'h5; //< 
    18'h13863: Data = 4'h2; //+ 
    18'h13864: Data = 4'h4; //> 
    18'h13865: Data = 4'h4; //> 
    18'h13866: Data = 4'h4; //> 
    18'h13867: Data = 4'h4; //> 
    18'h13868: Data = 4'h7; //] 
    18'h13869: Data = 4'h5; //< 
    18'h13870: Data = 4'h5; //< 
    18'h13871: Data = 4'h5; //< 
    18'h13872: Data = 4'h5; //< 
    18'h13873: Data = 4'h6; //[ 
    18'h13874: Data = 4'h3; //- 
    18'h13875: Data = 4'h4; //> 
    18'h13876: Data = 4'h4; //> 
    18'h13877: Data = 4'h4; //> 
    18'h13878: Data = 4'h4; //> 
    18'h13879: Data = 4'h2; //+ 
    18'h13880: Data = 4'h4; //> 
    18'h13881: Data = 4'h4; //> 
    18'h13882: Data = 4'h4; //> 
    18'h13883: Data = 4'h4; //> 
    18'h13884: Data = 4'h4; //> 
    18'h13885: Data = 4'h6; //[ 
    18'h13886: Data = 4'h4; //> 
    18'h13887: Data = 4'h2; //+ 
    18'h13888: Data = 4'h4; //> 
    18'h13889: Data = 4'h4; //> 
    18'h13890: Data = 4'h6; //[ 
    18'h13891: Data = 4'h3; //- 
    18'h13892: Data = 4'h5; //< 
    18'h13893: Data = 4'h5; //< 
    18'h13894: Data = 4'h3; //- 
    18'h13895: Data = 4'h4; //> 
    18'h13896: Data = 4'h4; //> 
    18'h13897: Data = 4'h7; //] 
    18'h13898: Data = 4'h5; //< 
    18'h13899: Data = 4'h5; //< 
    18'h13900: Data = 4'h6; //[ 
    18'h13901: Data = 4'h3; //- 
    18'h13902: Data = 4'h4; //> 
    18'h13903: Data = 4'h4; //> 
    18'h13904: Data = 4'h2; //+ 
    18'h13905: Data = 4'h5; //< 
    18'h13906: Data = 4'h5; //< 
    18'h13907: Data = 4'h7; //] 
    18'h13908: Data = 4'h4; //> 
    18'h13909: Data = 4'h4; //> 
    18'h13910: Data = 4'h4; //> 
    18'h13911: Data = 4'h4; //> 
    18'h13912: Data = 4'h4; //> 
    18'h13913: Data = 4'h4; //> 
    18'h13914: Data = 4'h4; //> 
    18'h13915: Data = 4'h4; //> 
    18'h13916: Data = 4'h7; //] 
    18'h13917: Data = 4'h5; //< 
    18'h13918: Data = 4'h5; //< 
    18'h13919: Data = 4'h5; //< 
    18'h13920: Data = 4'h5; //< 
    18'h13921: Data = 4'h5; //< 
    18'h13922: Data = 4'h5; //< 
    18'h13923: Data = 4'h5; //< 
    18'h13924: Data = 4'h5; //< 
    18'h13925: Data = 4'h2; //+ 
    18'h13926: Data = 4'h5; //< 
    18'h13927: Data = 4'h6; //[ 
    18'h13928: Data = 4'h4; //> 
    18'h13929: Data = 4'h6; //[ 
    18'h13930: Data = 4'h3; //- 
    18'h13931: Data = 4'h4; //> 
    18'h13932: Data = 4'h4; //> 
    18'h13933: Data = 4'h4; //> 
    18'h13934: Data = 4'h4; //> 
    18'h13935: Data = 4'h4; //> 
    18'h13936: Data = 4'h2; //+ 
    18'h13937: Data = 4'h5; //< 
    18'h13938: Data = 4'h5; //< 
    18'h13939: Data = 4'h5; //< 
    18'h13940: Data = 4'h5; //< 
    18'h13941: Data = 4'h6; //[ 
    18'h13942: Data = 4'h3; //- 
    18'h13943: Data = 4'h4; //> 
    18'h13944: Data = 4'h4; //> 
    18'h13945: Data = 4'h4; //> 
    18'h13946: Data = 4'h4; //> 
    18'h13947: Data = 4'h3; //- 
    18'h13948: Data = 4'h5; //< 
    18'h13949: Data = 4'h5; //< 
    18'h13950: Data = 4'h5; //< 
    18'h13951: Data = 4'h5; //< 
    18'h13952: Data = 4'h5; //< 
    18'h13953: Data = 4'h5; //< 
    18'h13954: Data = 4'h5; //< 
    18'h13955: Data = 4'h5; //< 
    18'h13956: Data = 4'h5; //< 
    18'h13957: Data = 4'h5; //< 
    18'h13958: Data = 4'h5; //< 
    18'h13959: Data = 4'h5; //< 
    18'h13960: Data = 4'h5; //< 
    18'h13961: Data = 4'h5; //< 
    18'h13962: Data = 4'h2; //+ 
    18'h13963: Data = 4'h4; //> 
    18'h13964: Data = 4'h4; //> 
    18'h13965: Data = 4'h4; //> 
    18'h13966: Data = 4'h4; //> 
    18'h13967: Data = 4'h4; //> 
    18'h13968: Data = 4'h4; //> 
    18'h13969: Data = 4'h4; //> 
    18'h13970: Data = 4'h4; //> 
    18'h13971: Data = 4'h4; //> 
    18'h13972: Data = 4'h4; //> 
    18'h13973: Data = 4'h4; //> 
    18'h13974: Data = 4'h6; //[ 
    18'h13975: Data = 4'h3; //- 
    18'h13976: Data = 4'h4; //> 
    18'h13977: Data = 4'h4; //> 
    18'h13978: Data = 4'h4; //> 
    18'h13979: Data = 4'h2; //+ 
    18'h13980: Data = 4'h5; //< 
    18'h13981: Data = 4'h5; //< 
    18'h13982: Data = 4'h5; //< 
    18'h13983: Data = 4'h7; //] 
    18'h13984: Data = 4'h5; //< 
    18'h13985: Data = 4'h7; //] 
    18'h13986: Data = 4'h4; //> 
    18'h13987: Data = 4'h6; //[ 
    18'h13988: Data = 4'h3; //- 
    18'h13989: Data = 4'h4; //> 
    18'h13990: Data = 4'h4; //> 
    18'h13991: Data = 4'h4; //> 
    18'h13992: Data = 4'h3; //- 
    18'h13993: Data = 4'h5; //< 
    18'h13994: Data = 4'h5; //< 
    18'h13995: Data = 4'h5; //< 
    18'h13996: Data = 4'h5; //< 
    18'h13997: Data = 4'h5; //< 
    18'h13998: Data = 4'h5; //< 
    18'h13999: Data = 4'h5; //< 
    18'h14000: Data = 4'h5; //< 
    18'h14001: Data = 4'h5; //< 
    18'h14002: Data = 4'h5; //< 
    18'h14003: Data = 4'h5; //< 
    18'h14004: Data = 4'h5; //< 
    18'h14005: Data = 4'h5; //< 
    18'h14006: Data = 4'h5; //< 
    18'h14007: Data = 4'h2; //+ 
    18'h14008: Data = 4'h4; //> 
    18'h14009: Data = 4'h4; //> 
    18'h14010: Data = 4'h4; //> 
    18'h14011: Data = 4'h4; //> 
    18'h14012: Data = 4'h4; //> 
    18'h14013: Data = 4'h4; //> 
    18'h14014: Data = 4'h4; //> 
    18'h14015: Data = 4'h4; //> 
    18'h14016: Data = 4'h4; //> 
    18'h14017: Data = 4'h4; //> 
    18'h14018: Data = 4'h4; //> 
    18'h14019: Data = 4'h7; //] 
    18'h14020: Data = 4'h5; //< 
    18'h14021: Data = 4'h5; //< 
    18'h14022: Data = 4'h7; //] 
    18'h14023: Data = 4'h4; //> 
    18'h14024: Data = 4'h6; //[ 
    18'h14025: Data = 4'h3; //- 
    18'h14026: Data = 4'h4; //> 
    18'h14027: Data = 4'h4; //> 
    18'h14028: Data = 4'h4; //> 
    18'h14029: Data = 4'h4; //> 
    18'h14030: Data = 4'h2; //+ 
    18'h14031: Data = 4'h5; //< 
    18'h14032: Data = 4'h5; //< 
    18'h14033: Data = 4'h5; //< 
    18'h14034: Data = 4'h6; //[ 
    18'h14035: Data = 4'h3; //- 
    18'h14036: Data = 4'h4; //> 
    18'h14037: Data = 4'h4; //> 
    18'h14038: Data = 4'h4; //> 
    18'h14039: Data = 4'h3; //- 
    18'h14040: Data = 4'h5; //< 
    18'h14041: Data = 4'h5; //< 
    18'h14042: Data = 4'h5; //< 
    18'h14043: Data = 4'h5; //< 
    18'h14044: Data = 4'h5; //< 
    18'h14045: Data = 4'h5; //< 
    18'h14046: Data = 4'h5; //< 
    18'h14047: Data = 4'h5; //< 
    18'h14048: Data = 4'h5; //< 
    18'h14049: Data = 4'h5; //< 
    18'h14050: Data = 4'h5; //< 
    18'h14051: Data = 4'h5; //< 
    18'h14052: Data = 4'h5; //< 
    18'h14053: Data = 4'h5; //< 
    18'h14054: Data = 4'h2; //+ 
    18'h14055: Data = 4'h4; //> 
    18'h14056: Data = 4'h4; //> 
    18'h14057: Data = 4'h4; //> 
    18'h14058: Data = 4'h4; //> 
    18'h14059: Data = 4'h4; //> 
    18'h14060: Data = 4'h4; //> 
    18'h14061: Data = 4'h4; //> 
    18'h14062: Data = 4'h4; //> 
    18'h14063: Data = 4'h4; //> 
    18'h14064: Data = 4'h4; //> 
    18'h14065: Data = 4'h4; //> 
    18'h14066: Data = 4'h7; //] 
    18'h14067: Data = 4'h5; //< 
    18'h14068: Data = 4'h7; //] 
    18'h14069: Data = 4'h4; //> 
    18'h14070: Data = 4'h6; //[ 
    18'h14071: Data = 4'h3; //- 
    18'h14072: Data = 4'h4; //> 
    18'h14073: Data = 4'h4; //> 
    18'h14074: Data = 4'h4; //> 
    18'h14075: Data = 4'h2; //+ 
    18'h14076: Data = 4'h5; //< 
    18'h14077: Data = 4'h5; //< 
    18'h14078: Data = 4'h5; //< 
    18'h14079: Data = 4'h7; //] 
    18'h14080: Data = 4'h5; //< 
    18'h14081: Data = 4'h5; //< 
    18'h14082: Data = 4'h5; //< 
    18'h14083: Data = 4'h5; //< 
    18'h14084: Data = 4'h5; //< 
    18'h14085: Data = 4'h5; //< 
    18'h14086: Data = 4'h5; //< 
    18'h14087: Data = 4'h5; //< 
    18'h14088: Data = 4'h5; //< 
    18'h14089: Data = 4'h5; //< 
    18'h14090: Data = 4'h5; //< 
    18'h14091: Data = 4'h5; //< 
    18'h14092: Data = 4'h7; //] 
    18'h14093: Data = 4'h4; //> 
    18'h14094: Data = 4'h4; //> 
    18'h14095: Data = 4'h4; //> 
    18'h14096: Data = 4'h4; //> 
    18'h14097: Data = 4'ha; //0 
    18'h14098: Data = 4'h5; //< 
    18'h14099: Data = 4'h5; //< 
    18'h14100: Data = 4'h5; //< 
    18'h14101: Data = 4'h5; //< 
    18'h14102: Data = 4'h7; //] 
    18'h14103: Data = 4'h4; //> 
    18'h14104: Data = 4'h4; //> 
    18'h14105: Data = 4'h4; //> 
    18'h14106: Data = 4'h6; //[ 
    18'h14107: Data = 4'h3; //- 
    18'h14108: Data = 4'h5; //< 
    18'h14109: Data = 4'h5; //< 
    18'h14110: Data = 4'h5; //< 
    18'h14111: Data = 4'h2; //+ 
    18'h14112: Data = 4'h4; //> 
    18'h14113: Data = 4'h4; //> 
    18'h14114: Data = 4'h4; //> 
    18'h14115: Data = 4'h7; //] 
    18'h14116: Data = 4'h5; //< 
    18'h14117: Data = 4'h5; //< 
    18'h14118: Data = 4'h5; //< 
    18'h14119: Data = 4'h6; //[ 
    18'h14120: Data = 4'h3; //- 
    18'h14121: Data = 4'h4; //> 
    18'h14122: Data = 4'h4; //> 
    18'h14123: Data = 4'h4; //> 
    18'h14124: Data = 4'h2; //+ 
    18'h14125: Data = 4'h4; //> 
    18'h14126: Data = 4'h4; //> 
    18'h14127: Data = 4'h4; //> 
    18'h14128: Data = 4'h4; //> 
    18'h14129: Data = 4'h4; //> 
    18'h14130: Data = 4'h4; //> 
    18'h14131: Data = 4'h6; //[ 
    18'h14132: Data = 4'h4; //> 
    18'h14133: Data = 4'h2; //+ 
    18'h14134: Data = 4'h4; //> 
    18'h14135: Data = 4'h6; //[ 
    18'h14136: Data = 4'h3; //- 
    18'h14137: Data = 4'h5; //< 
    18'h14138: Data = 4'h3; //- 
    18'h14139: Data = 4'h4; //> 
    18'h14140: Data = 4'h7; //] 
    18'h14141: Data = 4'h5; //< 
    18'h14142: Data = 4'h6; //[ 
    18'h14143: Data = 4'h3; //- 
    18'h14144: Data = 4'h4; //> 
    18'h14145: Data = 4'h2; //+ 
    18'h14146: Data = 4'h5; //< 
    18'h14147: Data = 4'h7; //] 
    18'h14148: Data = 4'h4; //> 
    18'h14149: Data = 4'h4; //> 
    18'h14150: Data = 4'h4; //> 
    18'h14151: Data = 4'h4; //> 
    18'h14152: Data = 4'h4; //> 
    18'h14153: Data = 4'h4; //> 
    18'h14154: Data = 4'h4; //> 
    18'h14155: Data = 4'h4; //> 
    18'h14156: Data = 4'h7; //] 
    18'h14157: Data = 4'h5; //< 
    18'h14158: Data = 4'h5; //< 
    18'h14159: Data = 4'h5; //< 
    18'h14160: Data = 4'h5; //< 
    18'h14161: Data = 4'h5; //< 
    18'h14162: Data = 4'h5; //< 
    18'h14163: Data = 4'h5; //< 
    18'h14164: Data = 4'h5; //< 
    18'h14165: Data = 4'h2; //+ 
    18'h14166: Data = 4'h5; //< 
    18'h14167: Data = 4'h6; //[ 
    18'h14168: Data = 4'h4; //> 
    18'h14169: Data = 4'h6; //[ 
    18'h14170: Data = 4'h3; //- 
    18'h14171: Data = 4'h4; //> 
    18'h14172: Data = 4'h4; //> 
    18'h14173: Data = 4'h4; //> 
    18'h14174: Data = 4'h4; //> 
    18'h14175: Data = 4'h4; //> 
    18'h14176: Data = 4'h2; //+ 
    18'h14177: Data = 4'h5; //< 
    18'h14178: Data = 4'h5; //< 
    18'h14179: Data = 4'h5; //< 
    18'h14180: Data = 4'h6; //[ 
    18'h14181: Data = 4'h3; //- 
    18'h14182: Data = 4'h4; //> 
    18'h14183: Data = 4'h4; //> 
    18'h14184: Data = 4'h4; //> 
    18'h14185: Data = 4'h3; //- 
    18'h14186: Data = 4'h5; //< 
    18'h14187: Data = 4'h5; //< 
    18'h14188: Data = 4'h5; //< 
    18'h14189: Data = 4'h5; //< 
    18'h14190: Data = 4'h5; //< 
    18'h14191: Data = 4'h5; //< 
    18'h14192: Data = 4'h5; //< 
    18'h14193: Data = 4'h5; //< 
    18'h14194: Data = 4'h5; //< 
    18'h14195: Data = 4'h5; //< 
    18'h14196: Data = 4'h5; //< 
    18'h14197: Data = 4'h5; //< 
    18'h14198: Data = 4'h5; //< 
    18'h14199: Data = 4'h5; //< 
    18'h14200: Data = 4'h2; //+ 
    18'h14201: Data = 4'h4; //> 
    18'h14202: Data = 4'h4; //> 
    18'h14203: Data = 4'h4; //> 
    18'h14204: Data = 4'h4; //> 
    18'h14205: Data = 4'h4; //> 
    18'h14206: Data = 4'h4; //> 
    18'h14207: Data = 4'h4; //> 
    18'h14208: Data = 4'h4; //> 
    18'h14209: Data = 4'h4; //> 
    18'h14210: Data = 4'h4; //> 
    18'h14211: Data = 4'h6; //[ 
    18'h14212: Data = 4'h3; //- 
    18'h14213: Data = 4'h4; //> 
    18'h14214: Data = 4'h4; //> 
    18'h14215: Data = 4'h4; //> 
    18'h14216: Data = 4'h4; //> 
    18'h14217: Data = 4'h2; //+ 
    18'h14218: Data = 4'h5; //< 
    18'h14219: Data = 4'h5; //< 
    18'h14220: Data = 4'h5; //< 
    18'h14221: Data = 4'h5; //< 
    18'h14222: Data = 4'h7; //] 
    18'h14223: Data = 4'h4; //> 
    18'h14224: Data = 4'h7; //] 
    18'h14225: Data = 4'h5; //< 
    18'h14226: Data = 4'h6; //[ 
    18'h14227: Data = 4'h3; //- 
    18'h14228: Data = 4'h4; //> 
    18'h14229: Data = 4'h4; //> 
    18'h14230: Data = 4'h4; //> 
    18'h14231: Data = 4'h4; //> 
    18'h14232: Data = 4'h3; //- 
    18'h14233: Data = 4'h5; //< 
    18'h14234: Data = 4'h5; //< 
    18'h14235: Data = 4'h5; //< 
    18'h14236: Data = 4'h5; //< 
    18'h14237: Data = 4'h5; //< 
    18'h14238: Data = 4'h5; //< 
    18'h14239: Data = 4'h5; //< 
    18'h14240: Data = 4'h5; //< 
    18'h14241: Data = 4'h5; //< 
    18'h14242: Data = 4'h5; //< 
    18'h14243: Data = 4'h5; //< 
    18'h14244: Data = 4'h5; //< 
    18'h14245: Data = 4'h5; //< 
    18'h14246: Data = 4'h5; //< 
    18'h14247: Data = 4'h2; //+ 
    18'h14248: Data = 4'h4; //> 
    18'h14249: Data = 4'h4; //> 
    18'h14250: Data = 4'h4; //> 
    18'h14251: Data = 4'h4; //> 
    18'h14252: Data = 4'h4; //> 
    18'h14253: Data = 4'h4; //> 
    18'h14254: Data = 4'h4; //> 
    18'h14255: Data = 4'h4; //> 
    18'h14256: Data = 4'h4; //> 
    18'h14257: Data = 4'h4; //> 
    18'h14258: Data = 4'h7; //] 
    18'h14259: Data = 4'h5; //< 
    18'h14260: Data = 4'h7; //] 
    18'h14261: Data = 4'h4; //> 
    18'h14262: Data = 4'h4; //> 
    18'h14263: Data = 4'h6; //[ 
    18'h14264: Data = 4'h3; //- 
    18'h14265: Data = 4'h4; //> 
    18'h14266: Data = 4'h4; //> 
    18'h14267: Data = 4'h4; //> 
    18'h14268: Data = 4'h2; //+ 
    18'h14269: Data = 4'h5; //< 
    18'h14270: Data = 4'h5; //< 
    18'h14271: Data = 4'h5; //< 
    18'h14272: Data = 4'h5; //< 
    18'h14273: Data = 4'h6; //[ 
    18'h14274: Data = 4'h3; //- 
    18'h14275: Data = 4'h4; //> 
    18'h14276: Data = 4'h4; //> 
    18'h14277: Data = 4'h4; //> 
    18'h14278: Data = 4'h4; //> 
    18'h14279: Data = 4'h3; //- 
    18'h14280: Data = 4'h5; //< 
    18'h14281: Data = 4'h5; //< 
    18'h14282: Data = 4'h5; //< 
    18'h14283: Data = 4'h5; //< 
    18'h14284: Data = 4'h5; //< 
    18'h14285: Data = 4'h5; //< 
    18'h14286: Data = 4'h5; //< 
    18'h14287: Data = 4'h5; //< 
    18'h14288: Data = 4'h5; //< 
    18'h14289: Data = 4'h5; //< 
    18'h14290: Data = 4'h5; //< 
    18'h14291: Data = 4'h5; //< 
    18'h14292: Data = 4'h5; //< 
    18'h14293: Data = 4'h5; //< 
    18'h14294: Data = 4'h2; //+ 
    18'h14295: Data = 4'h4; //> 
    18'h14296: Data = 4'h4; //> 
    18'h14297: Data = 4'h4; //> 
    18'h14298: Data = 4'h4; //> 
    18'h14299: Data = 4'h4; //> 
    18'h14300: Data = 4'h4; //> 
    18'h14301: Data = 4'h4; //> 
    18'h14302: Data = 4'h4; //> 
    18'h14303: Data = 4'h4; //> 
    18'h14304: Data = 4'h4; //> 
    18'h14305: Data = 4'h7; //] 
    18'h14306: Data = 4'h4; //> 
    18'h14307: Data = 4'h7; //] 
    18'h14308: Data = 4'h5; //< 
    18'h14309: Data = 4'h6; //[ 
    18'h14310: Data = 4'h3; //- 
    18'h14311: Data = 4'h4; //> 
    18'h14312: Data = 4'h4; //> 
    18'h14313: Data = 4'h4; //> 
    18'h14314: Data = 4'h4; //> 
    18'h14315: Data = 4'h2; //+ 
    18'h14316: Data = 4'h5; //< 
    18'h14317: Data = 4'h5; //< 
    18'h14318: Data = 4'h5; //< 
    18'h14319: Data = 4'h5; //< 
    18'h14320: Data = 4'h7; //] 
    18'h14321: Data = 4'h5; //< 
    18'h14322: Data = 4'h5; //< 
    18'h14323: Data = 4'h5; //< 
    18'h14324: Data = 4'h5; //< 
    18'h14325: Data = 4'h5; //< 
    18'h14326: Data = 4'h5; //< 
    18'h14327: Data = 4'h5; //< 
    18'h14328: Data = 4'h5; //< 
    18'h14329: Data = 4'h5; //< 
    18'h14330: Data = 4'h5; //< 
    18'h14331: Data = 4'h5; //< 
    18'h14332: Data = 4'h7; //] 
    18'h14333: Data = 4'h4; //> 
    18'h14334: Data = 4'h4; //> 
    18'h14335: Data = 4'h4; //> 
    18'h14336: Data = 4'h4; //> 
    18'h14337: Data = 4'h4; //> 
    18'h14338: Data = 4'h4; //> 
    18'h14339: Data = 4'h2; //+ 
    18'h14340: Data = 4'h5; //< 
    18'h14341: Data = 4'h5; //< 
    18'h14342: Data = 4'h5; //< 
    18'h14343: Data = 4'h5; //< 
    18'h14344: Data = 4'h5; //< 
    18'h14345: Data = 4'h5; //< 
    18'h14346: Data = 4'h7; //] 
    18'h14347: Data = 4'h7; //] 
    18'h14348: Data = 4'h4; //> 
    18'h14349: Data = 4'h4; //> 
    18'h14350: Data = 4'h4; //> 
    18'h14351: Data = 4'h4; //> 
    18'h14352: Data = 4'h6; //[ 
    18'h14353: Data = 4'h3; //- 
    18'h14354: Data = 4'h5; //< 
    18'h14355: Data = 4'h5; //< 
    18'h14356: Data = 4'h5; //< 
    18'h14357: Data = 4'h5; //< 
    18'h14358: Data = 4'h2; //+ 
    18'h14359: Data = 4'h4; //> 
    18'h14360: Data = 4'h4; //> 
    18'h14361: Data = 4'h4; //> 
    18'h14362: Data = 4'h4; //> 
    18'h14363: Data = 4'h7; //] 
    18'h14364: Data = 4'h5; //< 
    18'h14365: Data = 4'h5; //< 
    18'h14366: Data = 4'h5; //< 
    18'h14367: Data = 4'h5; //< 
    18'h14368: Data = 4'h6; //[ 
    18'h14369: Data = 4'h3; //- 
    18'h14370: Data = 4'h4; //> 
    18'h14371: Data = 4'h4; //> 
    18'h14372: Data = 4'h4; //> 
    18'h14373: Data = 4'h4; //> 
    18'h14374: Data = 4'h2; //+ 
    18'h14375: Data = 4'h4; //> 
    18'h14376: Data = 4'h4; //> 
    18'h14377: Data = 4'h4; //> 
    18'h14378: Data = 4'h4; //> 
    18'h14379: Data = 4'h4; //> 
    18'h14380: Data = 4'h6; //[ 
    18'h14381: Data = 4'h4; //> 
    18'h14382: Data = 4'h4; //> 
    18'h14383: Data = 4'h4; //> 
    18'h14384: Data = 4'h4; //> 
    18'h14385: Data = 4'h4; //> 
    18'h14386: Data = 4'h4; //> 
    18'h14387: Data = 4'h4; //> 
    18'h14388: Data = 4'h4; //> 
    18'h14389: Data = 4'h4; //> 
    18'h14390: Data = 4'h7; //] 
    18'h14391: Data = 4'h5; //< 
    18'h14392: Data = 4'h5; //< 
    18'h14393: Data = 4'h5; //< 
    18'h14394: Data = 4'h5; //< 
    18'h14395: Data = 4'h5; //< 
    18'h14396: Data = 4'h5; //< 
    18'h14397: Data = 4'h5; //< 
    18'h14398: Data = 4'h5; //< 
    18'h14399: Data = 4'h5; //< 
    18'h14400: Data = 4'h6; //[ 
    18'h14401: Data = 4'h4; //> 
    18'h14402: Data = 4'h6; //[ 
    18'h14403: Data = 4'h3; //- 
    18'h14404: Data = 4'h4; //> 
    18'h14405: Data = 4'h4; //> 
    18'h14406: Data = 4'h4; //> 
    18'h14407: Data = 4'h4; //> 
    18'h14408: Data = 4'h4; //> 
    18'h14409: Data = 4'h2; //+ 
    18'h14410: Data = 4'h5; //< 
    18'h14411: Data = 4'h5; //< 
    18'h14412: Data = 4'h5; //< 
    18'h14413: Data = 4'h5; //< 
    18'h14414: Data = 4'h6; //[ 
    18'h14415: Data = 4'h3; //- 
    18'h14416: Data = 4'h4; //> 
    18'h14417: Data = 4'h4; //> 
    18'h14418: Data = 4'h4; //> 
    18'h14419: Data = 4'h4; //> 
    18'h14420: Data = 4'h3; //- 
    18'h14421: Data = 4'h5; //< 
    18'h14422: Data = 4'h5; //< 
    18'h14423: Data = 4'h5; //< 
    18'h14424: Data = 4'h5; //< 
    18'h14425: Data = 4'h5; //< 
    18'h14426: Data = 4'h5; //< 
    18'h14427: Data = 4'h5; //< 
    18'h14428: Data = 4'h5; //< 
    18'h14429: Data = 4'h5; //< 
    18'h14430: Data = 4'h5; //< 
    18'h14431: Data = 4'h5; //< 
    18'h14432: Data = 4'h5; //< 
    18'h14433: Data = 4'h5; //< 
    18'h14434: Data = 4'h5; //< 
    18'h14435: Data = 4'h2; //+ 
    18'h14436: Data = 4'h4; //> 
    18'h14437: Data = 4'h4; //> 
    18'h14438: Data = 4'h4; //> 
    18'h14439: Data = 4'h4; //> 
    18'h14440: Data = 4'h4; //> 
    18'h14441: Data = 4'h4; //> 
    18'h14442: Data = 4'h4; //> 
    18'h14443: Data = 4'h4; //> 
    18'h14444: Data = 4'h4; //> 
    18'h14445: Data = 4'h4; //> 
    18'h14446: Data = 4'h4; //> 
    18'h14447: Data = 4'h6; //[ 
    18'h14448: Data = 4'h3; //- 
    18'h14449: Data = 4'h4; //> 
    18'h14450: Data = 4'h4; //> 
    18'h14451: Data = 4'h4; //> 
    18'h14452: Data = 4'h2; //+ 
    18'h14453: Data = 4'h5; //< 
    18'h14454: Data = 4'h5; //< 
    18'h14455: Data = 4'h5; //< 
    18'h14456: Data = 4'h7; //] 
    18'h14457: Data = 4'h5; //< 
    18'h14458: Data = 4'h7; //] 
    18'h14459: Data = 4'h4; //> 
    18'h14460: Data = 4'h6; //[ 
    18'h14461: Data = 4'h3; //- 
    18'h14462: Data = 4'h4; //> 
    18'h14463: Data = 4'h4; //> 
    18'h14464: Data = 4'h4; //> 
    18'h14465: Data = 4'h3; //- 
    18'h14466: Data = 4'h5; //< 
    18'h14467: Data = 4'h5; //< 
    18'h14468: Data = 4'h5; //< 
    18'h14469: Data = 4'h5; //< 
    18'h14470: Data = 4'h5; //< 
    18'h14471: Data = 4'h5; //< 
    18'h14472: Data = 4'h5; //< 
    18'h14473: Data = 4'h5; //< 
    18'h14474: Data = 4'h5; //< 
    18'h14475: Data = 4'h5; //< 
    18'h14476: Data = 4'h5; //< 
    18'h14477: Data = 4'h5; //< 
    18'h14478: Data = 4'h5; //< 
    18'h14479: Data = 4'h5; //< 
    18'h14480: Data = 4'h2; //+ 
    18'h14481: Data = 4'h4; //> 
    18'h14482: Data = 4'h4; //> 
    18'h14483: Data = 4'h4; //> 
    18'h14484: Data = 4'h4; //> 
    18'h14485: Data = 4'h4; //> 
    18'h14486: Data = 4'h4; //> 
    18'h14487: Data = 4'h4; //> 
    18'h14488: Data = 4'h4; //> 
    18'h14489: Data = 4'h4; //> 
    18'h14490: Data = 4'h4; //> 
    18'h14491: Data = 4'h4; //> 
    18'h14492: Data = 4'h7; //] 
    18'h14493: Data = 4'h5; //< 
    18'h14494: Data = 4'h5; //< 
    18'h14495: Data = 4'h7; //] 
    18'h14496: Data = 4'h4; //> 
    18'h14497: Data = 4'h6; //[ 
    18'h14498: Data = 4'h3; //- 
    18'h14499: Data = 4'h4; //> 
    18'h14500: Data = 4'h4; //> 
    18'h14501: Data = 4'h4; //> 
    18'h14502: Data = 4'h4; //> 
    18'h14503: Data = 4'h2; //+ 
    18'h14504: Data = 4'h5; //< 
    18'h14505: Data = 4'h5; //< 
    18'h14506: Data = 4'h5; //< 
    18'h14507: Data = 4'h6; //[ 
    18'h14508: Data = 4'h3; //- 
    18'h14509: Data = 4'h4; //> 
    18'h14510: Data = 4'h4; //> 
    18'h14511: Data = 4'h4; //> 
    18'h14512: Data = 4'h3; //- 
    18'h14513: Data = 4'h5; //< 
    18'h14514: Data = 4'h5; //< 
    18'h14515: Data = 4'h5; //< 
    18'h14516: Data = 4'h5; //< 
    18'h14517: Data = 4'h5; //< 
    18'h14518: Data = 4'h5; //< 
    18'h14519: Data = 4'h5; //< 
    18'h14520: Data = 4'h5; //< 
    18'h14521: Data = 4'h5; //< 
    18'h14522: Data = 4'h5; //< 
    18'h14523: Data = 4'h5; //< 
    18'h14524: Data = 4'h5; //< 
    18'h14525: Data = 4'h5; //< 
    18'h14526: Data = 4'h5; //< 
    18'h14527: Data = 4'h2; //+ 
    18'h14528: Data = 4'h4; //> 
    18'h14529: Data = 4'h4; //> 
    18'h14530: Data = 4'h4; //> 
    18'h14531: Data = 4'h4; //> 
    18'h14532: Data = 4'h4; //> 
    18'h14533: Data = 4'h4; //> 
    18'h14534: Data = 4'h4; //> 
    18'h14535: Data = 4'h4; //> 
    18'h14536: Data = 4'h4; //> 
    18'h14537: Data = 4'h4; //> 
    18'h14538: Data = 4'h4; //> 
    18'h14539: Data = 4'h7; //] 
    18'h14540: Data = 4'h5; //< 
    18'h14541: Data = 4'h7; //] 
    18'h14542: Data = 4'h4; //> 
    18'h14543: Data = 4'h6; //[ 
    18'h14544: Data = 4'h3; //- 
    18'h14545: Data = 4'h4; //> 
    18'h14546: Data = 4'h4; //> 
    18'h14547: Data = 4'h4; //> 
    18'h14548: Data = 4'h2; //+ 
    18'h14549: Data = 4'h5; //< 
    18'h14550: Data = 4'h5; //< 
    18'h14551: Data = 4'h5; //< 
    18'h14552: Data = 4'h7; //] 
    18'h14553: Data = 4'h5; //< 
    18'h14554: Data = 4'h5; //< 
    18'h14555: Data = 4'h5; //< 
    18'h14556: Data = 4'h5; //< 
    18'h14557: Data = 4'h5; //< 
    18'h14558: Data = 4'h5; //< 
    18'h14559: Data = 4'h5; //< 
    18'h14560: Data = 4'h5; //< 
    18'h14561: Data = 4'h5; //< 
    18'h14562: Data = 4'h5; //< 
    18'h14563: Data = 4'h5; //< 
    18'h14564: Data = 4'h5; //< 
    18'h14565: Data = 4'h7; //] 
    18'h14566: Data = 4'h7; //] 
    18'h14567: Data = 4'h4; //> 
    18'h14568: Data = 4'ha; //0 
    18'h14569: Data = 4'h4; //> 
    18'h14570: Data = 4'h4; //> 
    18'h14571: Data = 4'ha; //0 
    18'h14572: Data = 4'h4; //> 
    18'h14573: Data = 4'ha; //0 
    18'h14574: Data = 4'h4; //> 
    18'h14575: Data = 4'h4; //> 
    18'h14576: Data = 4'h4; //> 
    18'h14577: Data = 4'h4; //> 
    18'h14578: Data = 4'h4; //> 
    18'h14579: Data = 4'h6; //[ 
    18'h14580: Data = 4'h4; //> 
    18'h14581: Data = 4'h4; //> 
    18'h14582: Data = 4'ha; //0 
    18'h14583: Data = 4'h4; //> 
    18'h14584: Data = 4'ha; //0 
    18'h14585: Data = 4'h4; //> 
    18'h14586: Data = 4'h4; //> 
    18'h14587: Data = 4'h4; //> 
    18'h14588: Data = 4'h4; //> 
    18'h14589: Data = 4'h4; //> 
    18'h14590: Data = 4'h4; //> 
    18'h14591: Data = 4'h7; //] 
    18'h14592: Data = 4'h5; //< 
    18'h14593: Data = 4'h5; //< 
    18'h14594: Data = 4'h5; //< 
    18'h14595: Data = 4'h5; //< 
    18'h14596: Data = 4'h5; //< 
    18'h14597: Data = 4'h5; //< 
    18'h14598: Data = 4'h5; //< 
    18'h14599: Data = 4'h5; //< 
    18'h14600: Data = 4'h5; //< 
    18'h14601: Data = 4'h6; //[ 
    18'h14602: Data = 4'h5; //< 
    18'h14603: Data = 4'h5; //< 
    18'h14604: Data = 4'h5; //< 
    18'h14605: Data = 4'h5; //< 
    18'h14606: Data = 4'h5; //< 
    18'h14607: Data = 4'h5; //< 
    18'h14608: Data = 4'h5; //< 
    18'h14609: Data = 4'h5; //< 
    18'h14610: Data = 4'h5; //< 
    18'h14611: Data = 4'h7; //] 
    18'h14612: Data = 4'h4; //> 
    18'h14613: Data = 4'h4; //> 
    18'h14614: Data = 4'h4; //> 
    18'h14615: Data = 4'h4; //> 
    18'h14616: Data = 4'h4; //> 
    18'h14617: Data = 4'h4; //> 
    18'h14618: Data = 4'h4; //> 
    18'h14619: Data = 4'h4; //> 
    18'h14620: Data = 4'h4; //> 
    18'h14621: Data = 4'h6; //[ 
    18'h14622: Data = 4'h4; //> 
    18'h14623: Data = 4'h4; //> 
    18'h14624: Data = 4'h4; //> 
    18'h14625: Data = 4'h4; //> 
    18'h14626: Data = 4'h4; //> 
    18'h14627: Data = 4'h6; //[ 
    18'h14628: Data = 4'h3; //- 
    18'h14629: Data = 4'h5; //< 
    18'h14630: Data = 4'h5; //< 
    18'h14631: Data = 4'h5; //< 
    18'h14632: Data = 4'h5; //< 
    18'h14633: Data = 4'h2; //+ 
    18'h14634: Data = 4'h4; //> 
    18'h14635: Data = 4'h4; //> 
    18'h14636: Data = 4'h4; //> 
    18'h14637: Data = 4'h4; //> 
    18'h14638: Data = 4'h7; //] 
    18'h14639: Data = 4'h5; //< 
    18'h14640: Data = 4'h5; //< 
    18'h14641: Data = 4'h5; //< 
    18'h14642: Data = 4'h5; //< 
    18'h14643: Data = 4'h6; //[ 
    18'h14644: Data = 4'h3; //- 
    18'h14645: Data = 4'h4; //> 
    18'h14646: Data = 4'h4; //> 
    18'h14647: Data = 4'h4; //> 
    18'h14648: Data = 4'h4; //> 
    18'h14649: Data = 4'h2; //+ 
    18'h14650: Data = 4'h5; //< 
    18'h14651: Data = 4'h5; //< 
    18'h14652: Data = 4'h5; //< 
    18'h14653: Data = 4'h2; //+ 
    18'h14654: Data = 4'h5; //< 
    18'h14655: Data = 4'h7; //] 
    18'h14656: Data = 4'h4; //> 
    18'h14657: Data = 4'h4; //> 
    18'h14658: Data = 4'h4; //> 
    18'h14659: Data = 4'h4; //> 
    18'h14660: Data = 4'h4; //> 
    18'h14661: Data = 4'h4; //> 
    18'h14662: Data = 4'h4; //> 
    18'h14663: Data = 4'h4; //> 
    18'h14664: Data = 4'h7; //] 
    18'h14665: Data = 4'h5; //< 
    18'h14666: Data = 4'h5; //< 
    18'h14667: Data = 4'h5; //< 
    18'h14668: Data = 4'h5; //< 
    18'h14669: Data = 4'h5; //< 
    18'h14670: Data = 4'h5; //< 
    18'h14671: Data = 4'h5; //< 
    18'h14672: Data = 4'h5; //< 
    18'h14673: Data = 4'h5; //< 
    18'h14674: Data = 4'h6; //[ 
    18'h14675: Data = 4'h5; //< 
    18'h14676: Data = 4'h5; //< 
    18'h14677: Data = 4'h5; //< 
    18'h14678: Data = 4'h5; //< 
    18'h14679: Data = 4'h5; //< 
    18'h14680: Data = 4'h5; //< 
    18'h14681: Data = 4'h5; //< 
    18'h14682: Data = 4'h5; //< 
    18'h14683: Data = 4'h5; //< 
    18'h14684: Data = 4'h7; //] 
    18'h14685: Data = 4'h4; //> 
    18'h14686: Data = 4'h4; //> 
    18'h14687: Data = 4'h4; //> 
    18'h14688: Data = 4'h4; //> 
    18'h14689: Data = 4'h4; //> 
    18'h14690: Data = 4'h4; //> 
    18'h14691: Data = 4'h4; //> 
    18'h14692: Data = 4'h4; //> 
    18'h14693: Data = 4'h4; //> 
    18'h14694: Data = 4'h2; //+ 
    18'h14695: Data = 4'h2; //+ 
    18'h14696: Data = 4'h2; //+ 
    18'h14697: Data = 4'h2; //+ 
    18'h14698: Data = 4'h2; //+ 
    18'h14699: Data = 4'h2; //+ 
    18'h14700: Data = 4'h2; //+ 
    18'h14701: Data = 4'h2; //+ 
    18'h14702: Data = 4'h2; //+ 
    18'h14703: Data = 4'h2; //+ 
    18'h14704: Data = 4'h2; //+ 
    18'h14705: Data = 4'h2; //+ 
    18'h14706: Data = 4'h2; //+ 
    18'h14707: Data = 4'h2; //+ 
    18'h14708: Data = 4'h2; //+ 
    18'h14709: Data = 4'h6; //[ 
    18'h14710: Data = 4'h6; //[ 
    18'h14711: Data = 4'h4; //> 
    18'h14712: Data = 4'h4; //> 
    18'h14713: Data = 4'h4; //> 
    18'h14714: Data = 4'h4; //> 
    18'h14715: Data = 4'h4; //> 
    18'h14716: Data = 4'h4; //> 
    18'h14717: Data = 4'h4; //> 
    18'h14718: Data = 4'h4; //> 
    18'h14719: Data = 4'h4; //> 
    18'h14720: Data = 4'h7; //] 
    18'h14721: Data = 4'h2; //+ 
    18'h14722: Data = 4'h4; //> 
    18'h14723: Data = 4'ha; //0 
    18'h14724: Data = 4'h4; //> 
    18'h14725: Data = 4'ha; //0 
    18'h14726: Data = 4'h4; //> 
    18'h14727: Data = 4'ha; //0 
    18'h14728: Data = 4'h4; //> 
    18'h14729: Data = 4'ha; //0 
    18'h14730: Data = 4'h4; //> 
    18'h14731: Data = 4'ha; //0 
    18'h14732: Data = 4'h4; //> 
    18'h14733: Data = 4'ha; //0 
    18'h14734: Data = 4'h4; //> 
    18'h14735: Data = 4'ha; //0 
    18'h14736: Data = 4'h4; //> 
    18'h14737: Data = 4'ha; //0 
    18'h14738: Data = 4'h4; //> 
    18'h14739: Data = 4'ha; //0 
    18'h14740: Data = 4'h5; //< 
    18'h14741: Data = 4'h5; //< 
    18'h14742: Data = 4'h5; //< 
    18'h14743: Data = 4'h5; //< 
    18'h14744: Data = 4'h5; //< 
    18'h14745: Data = 4'h5; //< 
    18'h14746: Data = 4'h5; //< 
    18'h14747: Data = 4'h5; //< 
    18'h14748: Data = 4'h5; //< 
    18'h14749: Data = 4'h6; //[ 
    18'h14750: Data = 4'h5; //< 
    18'h14751: Data = 4'h5; //< 
    18'h14752: Data = 4'h5; //< 
    18'h14753: Data = 4'h5; //< 
    18'h14754: Data = 4'h5; //< 
    18'h14755: Data = 4'h5; //< 
    18'h14756: Data = 4'h5; //< 
    18'h14757: Data = 4'h5; //< 
    18'h14758: Data = 4'h5; //< 
    18'h14759: Data = 4'h7; //] 
    18'h14760: Data = 4'h4; //> 
    18'h14761: Data = 4'h4; //> 
    18'h14762: Data = 4'h4; //> 
    18'h14763: Data = 4'h4; //> 
    18'h14764: Data = 4'h4; //> 
    18'h14765: Data = 4'h4; //> 
    18'h14766: Data = 4'h4; //> 
    18'h14767: Data = 4'h4; //> 
    18'h14768: Data = 4'h4; //> 
    18'h14769: Data = 4'h3; //- 
    18'h14770: Data = 4'h7; //] 
    18'h14771: Data = 4'h2; //+ 
    18'h14772: Data = 4'h6; //[ 
    18'h14773: Data = 4'h4; //> 
    18'h14774: Data = 4'h2; //+ 
    18'h14775: Data = 4'h4; //> 
    18'h14776: Data = 4'h4; //> 
    18'h14777: Data = 4'h4; //> 
    18'h14778: Data = 4'h4; //> 
    18'h14779: Data = 4'h4; //> 
    18'h14780: Data = 4'h4; //> 
    18'h14781: Data = 4'h4; //> 
    18'h14782: Data = 4'h4; //> 
    18'h14783: Data = 4'h7; //] 
    18'h14784: Data = 4'h5; //< 
    18'h14785: Data = 4'h5; //< 
    18'h14786: Data = 4'h5; //< 
    18'h14787: Data = 4'h5; //< 
    18'h14788: Data = 4'h5; //< 
    18'h14789: Data = 4'h5; //< 
    18'h14790: Data = 4'h5; //< 
    18'h14791: Data = 4'h5; //< 
    18'h14792: Data = 4'h5; //< 
    18'h14793: Data = 4'h6; //[ 
    18'h14794: Data = 4'h5; //< 
    18'h14795: Data = 4'h5; //< 
    18'h14796: Data = 4'h5; //< 
    18'h14797: Data = 4'h5; //< 
    18'h14798: Data = 4'h5; //< 
    18'h14799: Data = 4'h5; //< 
    18'h14800: Data = 4'h5; //< 
    18'h14801: Data = 4'h5; //< 
    18'h14802: Data = 4'h5; //< 
    18'h14803: Data = 4'h7; //] 
    18'h14804: Data = 4'h4; //> 
    18'h14805: Data = 4'h4; //> 
    18'h14806: Data = 4'h4; //> 
    18'h14807: Data = 4'h4; //> 
    18'h14808: Data = 4'h4; //> 
    18'h14809: Data = 4'h4; //> 
    18'h14810: Data = 4'h4; //> 
    18'h14811: Data = 4'h4; //> 
    18'h14812: Data = 4'h4; //> 
    18'h14813: Data = 4'h6; //[ 
    18'h14814: Data = 4'h4; //> 
    18'h14815: Data = 4'h3; //- 
    18'h14816: Data = 4'h4; //> 
    18'h14817: Data = 4'h4; //> 
    18'h14818: Data = 4'h4; //> 
    18'h14819: Data = 4'h4; //> 
    18'h14820: Data = 4'h6; //[ 
    18'h14821: Data = 4'h3; //- 
    18'h14822: Data = 4'h5; //< 
    18'h14823: Data = 4'h5; //< 
    18'h14824: Data = 4'h5; //< 
    18'h14825: Data = 4'h5; //< 
    18'h14826: Data = 4'h2; //+ 
    18'h14827: Data = 4'h4; //> 
    18'h14828: Data = 4'h4; //> 
    18'h14829: Data = 4'h4; //> 
    18'h14830: Data = 4'h4; //> 
    18'h14831: Data = 4'h7; //] 
    18'h14832: Data = 4'h5; //< 
    18'h14833: Data = 4'h5; //< 
    18'h14834: Data = 4'h5; //< 
    18'h14835: Data = 4'h5; //< 
    18'h14836: Data = 4'h6; //[ 
    18'h14837: Data = 4'h3; //- 
    18'h14838: Data = 4'h4; //> 
    18'h14839: Data = 4'h4; //> 
    18'h14840: Data = 4'h4; //> 
    18'h14841: Data = 4'h4; //> 
    18'h14842: Data = 4'h2; //+ 
    18'h14843: Data = 4'h5; //< 
    18'h14844: Data = 4'h5; //< 
    18'h14845: Data = 4'h5; //< 
    18'h14846: Data = 4'h5; //< 
    18'h14847: Data = 4'h5; //< 
    18'h14848: Data = 4'h6; //[ 
    18'h14849: Data = 4'h3; //- 
    18'h14850: Data = 4'h4; //> 
    18'h14851: Data = 4'h4; //> 
    18'h14852: Data = 4'h6; //[ 
    18'h14853: Data = 4'h3; //- 
    18'h14854: Data = 4'h5; //< 
    18'h14855: Data = 4'h5; //< 
    18'h14856: Data = 4'h2; //+ 
    18'h14857: Data = 4'h4; //> 
    18'h14858: Data = 4'h4; //> 
    18'h14859: Data = 4'h7; //] 
    18'h14860: Data = 4'h5; //< 
    18'h14861: Data = 4'h5; //< 
    18'h14862: Data = 4'h6; //[ 
    18'h14863: Data = 4'h3; //- 
    18'h14864: Data = 4'h4; //> 
    18'h14865: Data = 4'h4; //> 
    18'h14866: Data = 4'h2; //+ 
    18'h14867: Data = 4'h4; //> 
    18'h14868: Data = 4'h2; //+ 
    18'h14869: Data = 4'h5; //< 
    18'h14870: Data = 4'h5; //< 
    18'h14871: Data = 4'h5; //< 
    18'h14872: Data = 4'h7; //] 
    18'h14873: Data = 4'h2; //+ 
    18'h14874: Data = 4'h4; //> 
    18'h14875: Data = 4'h4; //> 
    18'h14876: Data = 4'h4; //> 
    18'h14877: Data = 4'h4; //> 
    18'h14878: Data = 4'h4; //> 
    18'h14879: Data = 4'h4; //> 
    18'h14880: Data = 4'h4; //> 
    18'h14881: Data = 4'h4; //> 
    18'h14882: Data = 4'h4; //> 
    18'h14883: Data = 4'h7; //] 
    18'h14884: Data = 4'h5; //< 
    18'h14885: Data = 4'h5; //< 
    18'h14886: Data = 4'h5; //< 
    18'h14887: Data = 4'h5; //< 
    18'h14888: Data = 4'h5; //< 
    18'h14889: Data = 4'h5; //< 
    18'h14890: Data = 4'h5; //< 
    18'h14891: Data = 4'h5; //< 
    18'h14892: Data = 4'h6; //[ 
    18'h14893: Data = 4'h5; //< 
    18'h14894: Data = 4'h5; //< 
    18'h14895: Data = 4'h5; //< 
    18'h14896: Data = 4'h5; //< 
    18'h14897: Data = 4'h5; //< 
    18'h14898: Data = 4'h5; //< 
    18'h14899: Data = 4'h5; //< 
    18'h14900: Data = 4'h5; //< 
    18'h14901: Data = 4'h5; //< 
    18'h14902: Data = 4'h7; //] 
    18'h14903: Data = 4'h7; //] 
    18'h14904: Data = 4'h4; //> 
    18'h14905: Data = 4'h4; //> 
    18'h14906: Data = 4'h4; //> 
    18'h14907: Data = 4'h4; //> 
    18'h14908: Data = 4'h4; //> 
    18'h14909: Data = 4'h4; //> 
    18'h14910: Data = 4'h4; //> 
    18'h14911: Data = 4'h4; //> 
    18'h14912: Data = 4'h4; //> 
    18'h14913: Data = 4'h6; //[ 
    18'h14914: Data = 4'h4; //> 
    18'h14915: Data = 4'h4; //> 
    18'h14916: Data = 4'h4; //> 
    18'h14917: Data = 4'h4; //> 
    18'h14918: Data = 4'h4; //> 
    18'h14919: Data = 4'h4; //> 
    18'h14920: Data = 4'h4; //> 
    18'h14921: Data = 4'h4; //> 
    18'h14922: Data = 4'h4; //> 
    18'h14923: Data = 4'h7; //] 
    18'h14924: Data = 4'h5; //< 
    18'h14925: Data = 4'h5; //< 
    18'h14926: Data = 4'h5; //< 
    18'h14927: Data = 4'h5; //< 
    18'h14928: Data = 4'h5; //< 
    18'h14929: Data = 4'h5; //< 
    18'h14930: Data = 4'h5; //< 
    18'h14931: Data = 4'h5; //< 
    18'h14932: Data = 4'h5; //< 
    18'h14933: Data = 4'h6; //[ 
    18'h14934: Data = 4'h4; //> 
    18'h14935: Data = 4'h6; //[ 
    18'h14936: Data = 4'h3; //- 
    18'h14937: Data = 4'h4; //> 
    18'h14938: Data = 4'h4; //> 
    18'h14939: Data = 4'h4; //> 
    18'h14940: Data = 4'h4; //> 
    18'h14941: Data = 4'h4; //> 
    18'h14942: Data = 4'h4; //> 
    18'h14943: Data = 4'h4; //> 
    18'h14944: Data = 4'h4; //> 
    18'h14945: Data = 4'h4; //> 
    18'h14946: Data = 4'h2; //+ 
    18'h14947: Data = 4'h5; //< 
    18'h14948: Data = 4'h5; //< 
    18'h14949: Data = 4'h5; //< 
    18'h14950: Data = 4'h5; //< 
    18'h14951: Data = 4'h5; //< 
    18'h14952: Data = 4'h5; //< 
    18'h14953: Data = 4'h5; //< 
    18'h14954: Data = 4'h5; //< 
    18'h14955: Data = 4'h5; //< 
    18'h14956: Data = 4'h7; //] 
    18'h14957: Data = 4'h5; //< 
    18'h14958: Data = 4'h5; //< 
    18'h14959: Data = 4'h5; //< 
    18'h14960: Data = 4'h5; //< 
    18'h14961: Data = 4'h5; //< 
    18'h14962: Data = 4'h5; //< 
    18'h14963: Data = 4'h5; //< 
    18'h14964: Data = 4'h5; //< 
    18'h14965: Data = 4'h5; //< 
    18'h14966: Data = 4'h5; //< 
    18'h14967: Data = 4'h7; //] 
    18'h14968: Data = 4'h4; //> 
    18'h14969: Data = 4'h6; //[ 
    18'h14970: Data = 4'h3; //- 
    18'h14971: Data = 4'h4; //> 
    18'h14972: Data = 4'h4; //> 
    18'h14973: Data = 4'h4; //> 
    18'h14974: Data = 4'h4; //> 
    18'h14975: Data = 4'h4; //> 
    18'h14976: Data = 4'h4; //> 
    18'h14977: Data = 4'h4; //> 
    18'h14978: Data = 4'h4; //> 
    18'h14979: Data = 4'h4; //> 
    18'h14980: Data = 4'h2; //+ 
    18'h14981: Data = 4'h5; //< 
    18'h14982: Data = 4'h5; //< 
    18'h14983: Data = 4'h5; //< 
    18'h14984: Data = 4'h5; //< 
    18'h14985: Data = 4'h5; //< 
    18'h14986: Data = 4'h5; //< 
    18'h14987: Data = 4'h5; //< 
    18'h14988: Data = 4'h5; //< 
    18'h14989: Data = 4'h5; //< 
    18'h14990: Data = 4'h7; //] 
    18'h14991: Data = 4'h5; //< 
    18'h14992: Data = 4'h2; //+ 
    18'h14993: Data = 4'h4; //> 
    18'h14994: Data = 4'h4; //> 
    18'h14995: Data = 4'h4; //> 
    18'h14996: Data = 4'h4; //> 
    18'h14997: Data = 4'h4; //> 
    18'h14998: Data = 4'h4; //> 
    18'h14999: Data = 4'h4; //> 
    18'h15000: Data = 4'h4; //> 
    18'h15001: Data = 4'h7; //] 
    18'h15002: Data = 4'h5; //< 
    18'h15003: Data = 4'h5; //< 
    18'h15004: Data = 4'h5; //< 
    18'h15005: Data = 4'h5; //< 
    18'h15006: Data = 4'h5; //< 
    18'h15007: Data = 4'h5; //< 
    18'h15008: Data = 4'h5; //< 
    18'h15009: Data = 4'h5; //< 
    18'h15010: Data = 4'h5; //< 
    18'h15011: Data = 4'h6; //[ 
    18'h15012: Data = 4'h4; //> 
    18'h15013: Data = 4'ha; //0 
    18'h15014: Data = 4'h5; //< 
    18'h15015: Data = 4'h3; //- 
    18'h15016: Data = 4'h4; //> 
    18'h15017: Data = 4'h4; //> 
    18'h15018: Data = 4'h4; //> 
    18'h15019: Data = 4'h6; //[ 
    18'h15020: Data = 4'h3; //- 
    18'h15021: Data = 4'h5; //< 
    18'h15022: Data = 4'h5; //< 
    18'h15023: Data = 4'h5; //< 
    18'h15024: Data = 4'h2; //+ 
    18'h15025: Data = 4'h4; //> 
    18'h15026: Data = 4'h6; //[ 
    18'h15027: Data = 4'h5; //< 
    18'h15028: Data = 4'h3; //- 
    18'h15029: Data = 4'h4; //> 
    18'h15030: Data = 4'h3; //- 
    18'h15031: Data = 4'h5; //< 
    18'h15032: Data = 4'h5; //< 
    18'h15033: Data = 4'h5; //< 
    18'h15034: Data = 4'h5; //< 
    18'h15035: Data = 4'h5; //< 
    18'h15036: Data = 4'h5; //< 
    18'h15037: Data = 4'h5; //< 
    18'h15038: Data = 4'h2; //+ 
    18'h15039: Data = 4'h4; //> 
    18'h15040: Data = 4'h4; //> 
    18'h15041: Data = 4'h4; //> 
    18'h15042: Data = 4'h4; //> 
    18'h15043: Data = 4'h4; //> 
    18'h15044: Data = 4'h4; //> 
    18'h15045: Data = 4'h4; //> 
    18'h15046: Data = 4'h7; //] 
    18'h15047: Data = 4'h5; //< 
    18'h15048: Data = 4'h6; //[ 
    18'h15049: Data = 4'h3; //- 
    18'h15050: Data = 4'h4; //> 
    18'h15051: Data = 4'h2; //+ 
    18'h15052: Data = 4'h5; //< 
    18'h15053: Data = 4'h7; //] 
    18'h15054: Data = 4'h4; //> 
    18'h15055: Data = 4'h4; //> 
    18'h15056: Data = 4'h4; //> 
    18'h15057: Data = 4'h7; //] 
    18'h15058: Data = 4'h5; //< 
    18'h15059: Data = 4'h5; //< 
    18'h15060: Data = 4'h6; //[ 
    18'h15061: Data = 4'h3; //- 
    18'h15062: Data = 4'h4; //> 
    18'h15063: Data = 4'h4; //> 
    18'h15064: Data = 4'h2; //+ 
    18'h15065: Data = 4'h5; //< 
    18'h15066: Data = 4'h5; //< 
    18'h15067: Data = 4'h7; //] 
    18'h15068: Data = 4'h5; //< 
    18'h15069: Data = 4'h2; //+ 
    18'h15070: Data = 4'h5; //< 
    18'h15071: Data = 4'h5; //< 
    18'h15072: Data = 4'h5; //< 
    18'h15073: Data = 4'h5; //< 
    18'h15074: Data = 4'h5; //< 
    18'h15075: Data = 4'h5; //< 
    18'h15076: Data = 4'h5; //< 
    18'h15077: Data = 4'h5; //< 
    18'h15078: Data = 4'h5; //< 
    18'h15079: Data = 4'h7; //] 
    18'h15080: Data = 4'h4; //> 
    18'h15081: Data = 4'h4; //> 
    18'h15082: Data = 4'h4; //> 
    18'h15083: Data = 4'h4; //> 
    18'h15084: Data = 4'h4; //> 
    18'h15085: Data = 4'h4; //> 
    18'h15086: Data = 4'h4; //> 
    18'h15087: Data = 4'h4; //> 
    18'h15088: Data = 4'h4; //> 
    18'h15089: Data = 4'h6; //[ 
    18'h15090: Data = 4'h4; //> 
    18'h15091: Data = 4'h4; //> 
    18'h15092: Data = 4'h4; //> 
    18'h15093: Data = 4'h6; //[ 
    18'h15094: Data = 4'h3; //- 
    18'h15095: Data = 4'h5; //< 
    18'h15096: Data = 4'h5; //< 
    18'h15097: Data = 4'h5; //< 
    18'h15098: Data = 4'h5; //< 
    18'h15099: Data = 4'h5; //< 
    18'h15100: Data = 4'h5; //< 
    18'h15101: Data = 4'h5; //< 
    18'h15102: Data = 4'h5; //< 
    18'h15103: Data = 4'h5; //< 
    18'h15104: Data = 4'h5; //< 
    18'h15105: Data = 4'h5; //< 
    18'h15106: Data = 4'h5; //< 
    18'h15107: Data = 4'h5; //< 
    18'h15108: Data = 4'h5; //< 
    18'h15109: Data = 4'h5; //< 
    18'h15110: Data = 4'h5; //< 
    18'h15111: Data = 4'h5; //< 
    18'h15112: Data = 4'h5; //< 
    18'h15113: Data = 4'h5; //< 
    18'h15114: Data = 4'h5; //< 
    18'h15115: Data = 4'h5; //< 
    18'h15116: Data = 4'h5; //< 
    18'h15117: Data = 4'h5; //< 
    18'h15118: Data = 4'h5; //< 
    18'h15119: Data = 4'h5; //< 
    18'h15120: Data = 4'h5; //< 
    18'h15121: Data = 4'h5; //< 
    18'h15122: Data = 4'h5; //< 
    18'h15123: Data = 4'h5; //< 
    18'h15124: Data = 4'h5; //< 
    18'h15125: Data = 4'h5; //< 
    18'h15126: Data = 4'h5; //< 
    18'h15127: Data = 4'h5; //< 
    18'h15128: Data = 4'h5; //< 
    18'h15129: Data = 4'h5; //< 
    18'h15130: Data = 4'h5; //< 
    18'h15131: Data = 4'h2; //+ 
    18'h15132: Data = 4'h4; //> 
    18'h15133: Data = 4'h4; //> 
    18'h15134: Data = 4'h4; //> 
    18'h15135: Data = 4'h4; //> 
    18'h15136: Data = 4'h4; //> 
    18'h15137: Data = 4'h4; //> 
    18'h15138: Data = 4'h4; //> 
    18'h15139: Data = 4'h4; //> 
    18'h15140: Data = 4'h4; //> 
    18'h15141: Data = 4'h4; //> 
    18'h15142: Data = 4'h4; //> 
    18'h15143: Data = 4'h4; //> 
    18'h15144: Data = 4'h4; //> 
    18'h15145: Data = 4'h4; //> 
    18'h15146: Data = 4'h4; //> 
    18'h15147: Data = 4'h4; //> 
    18'h15148: Data = 4'h4; //> 
    18'h15149: Data = 4'h4; //> 
    18'h15150: Data = 4'h4; //> 
    18'h15151: Data = 4'h4; //> 
    18'h15152: Data = 4'h4; //> 
    18'h15153: Data = 4'h4; //> 
    18'h15154: Data = 4'h4; //> 
    18'h15155: Data = 4'h4; //> 
    18'h15156: Data = 4'h4; //> 
    18'h15157: Data = 4'h4; //> 
    18'h15158: Data = 4'h4; //> 
    18'h15159: Data = 4'h4; //> 
    18'h15160: Data = 4'h4; //> 
    18'h15161: Data = 4'h4; //> 
    18'h15162: Data = 4'h4; //> 
    18'h15163: Data = 4'h4; //> 
    18'h15164: Data = 4'h4; //> 
    18'h15165: Data = 4'h4; //> 
    18'h15166: Data = 4'h4; //> 
    18'h15167: Data = 4'h4; //> 
    18'h15168: Data = 4'h7; //] 
    18'h15169: Data = 4'h4; //> 
    18'h15170: Data = 4'h4; //> 
    18'h15171: Data = 4'h4; //> 
    18'h15172: Data = 4'h4; //> 
    18'h15173: Data = 4'h4; //> 
    18'h15174: Data = 4'h4; //> 
    18'h15175: Data = 4'h7; //] 
    18'h15176: Data = 4'h5; //< 
    18'h15177: Data = 4'h5; //< 
    18'h15178: Data = 4'h5; //< 
    18'h15179: Data = 4'h5; //< 
    18'h15180: Data = 4'h5; //< 
    18'h15181: Data = 4'h5; //< 
    18'h15182: Data = 4'h5; //< 
    18'h15183: Data = 4'h5; //< 
    18'h15184: Data = 4'h5; //< 
    18'h15185: Data = 4'h6; //[ 
    18'h15186: Data = 4'h5; //< 
    18'h15187: Data = 4'h5; //< 
    18'h15188: Data = 4'h5; //< 
    18'h15189: Data = 4'h5; //< 
    18'h15190: Data = 4'h5; //< 
    18'h15191: Data = 4'h5; //< 
    18'h15192: Data = 4'h5; //< 
    18'h15193: Data = 4'h5; //< 
    18'h15194: Data = 4'h5; //< 
    18'h15195: Data = 4'h7; //] 
    18'h15196: Data = 4'h4; //> 
    18'h15197: Data = 4'h4; //> 
    18'h15198: Data = 4'h4; //> 
    18'h15199: Data = 4'h4; //> 
    18'h15200: Data = 4'h4; //> 
    18'h15201: Data = 4'ha; //0 
    18'h15202: Data = 4'h4; //> 
    18'h15203: Data = 4'h4; //> 
    18'h15204: Data = 4'h4; //> 
    18'h15205: Data = 4'h4; //> 
    18'h15206: Data = 4'h2; //+ 
    18'h15207: Data = 4'h2; //+ 
    18'h15208: Data = 4'h2; //+ 
    18'h15209: Data = 4'h2; //+ 
    18'h15210: Data = 4'h2; //+ 
    18'h15211: Data = 4'h2; //+ 
    18'h15212: Data = 4'h2; //+ 
    18'h15213: Data = 4'h2; //+ 
    18'h15214: Data = 4'h2; //+ 
    18'h15215: Data = 4'h2; //+ 
    18'h15216: Data = 4'h2; //+ 
    18'h15217: Data = 4'h2; //+ 
    18'h15218: Data = 4'h2; //+ 
    18'h15219: Data = 4'h2; //+ 
    18'h15220: Data = 4'h2; //+ 
    18'h15221: Data = 4'h6; //[ 
    18'h15222: Data = 4'h6; //[ 
    18'h15223: Data = 4'h4; //> 
    18'h15224: Data = 4'h4; //> 
    18'h15225: Data = 4'h4; //> 
    18'h15226: Data = 4'h4; //> 
    18'h15227: Data = 4'h4; //> 
    18'h15228: Data = 4'h4; //> 
    18'h15229: Data = 4'h4; //> 
    18'h15230: Data = 4'h4; //> 
    18'h15231: Data = 4'h4; //> 
    18'h15232: Data = 4'h7; //] 
    18'h15233: Data = 4'h5; //< 
    18'h15234: Data = 4'h5; //< 
    18'h15235: Data = 4'h5; //< 
    18'h15236: Data = 4'h5; //< 
    18'h15237: Data = 4'h5; //< 
    18'h15238: Data = 4'h5; //< 
    18'h15239: Data = 4'h5; //< 
    18'h15240: Data = 4'h5; //< 
    18'h15241: Data = 4'h5; //< 
    18'h15242: Data = 4'h3; //- 
    18'h15243: Data = 4'h5; //< 
    18'h15244: Data = 4'h5; //< 
    18'h15245: Data = 4'h5; //< 
    18'h15246: Data = 4'h5; //< 
    18'h15247: Data = 4'h5; //< 
    18'h15248: Data = 4'h5; //< 
    18'h15249: Data = 4'h5; //< 
    18'h15250: Data = 4'h5; //< 
    18'h15251: Data = 4'h5; //< 
    18'h15252: Data = 4'h6; //[ 
    18'h15253: Data = 4'h5; //< 
    18'h15254: Data = 4'h5; //< 
    18'h15255: Data = 4'h5; //< 
    18'h15256: Data = 4'h5; //< 
    18'h15257: Data = 4'h5; //< 
    18'h15258: Data = 4'h5; //< 
    18'h15259: Data = 4'h5; //< 
    18'h15260: Data = 4'h5; //< 
    18'h15261: Data = 4'h5; //< 
    18'h15262: Data = 4'h7; //] 
    18'h15263: Data = 4'h4; //> 
    18'h15264: Data = 4'h4; //> 
    18'h15265: Data = 4'h4; //> 
    18'h15266: Data = 4'h4; //> 
    18'h15267: Data = 4'h4; //> 
    18'h15268: Data = 4'h4; //> 
    18'h15269: Data = 4'h4; //> 
    18'h15270: Data = 4'h4; //> 
    18'h15271: Data = 4'h4; //> 
    18'h15272: Data = 4'h3; //- 
    18'h15273: Data = 4'h7; //] 
    18'h15274: Data = 4'h2; //+ 
    18'h15275: Data = 4'h6; //[ 
    18'h15276: Data = 4'h4; //> 
    18'h15277: Data = 4'h4; //> 
    18'h15278: Data = 4'h4; //> 
    18'h15279: Data = 4'h6; //[ 
    18'h15280: Data = 4'h3; //- 
    18'h15281: Data = 4'h5; //< 
    18'h15282: Data = 4'h5; //< 
    18'h15283: Data = 4'h5; //< 
    18'h15284: Data = 4'h3; //- 
    18'h15285: Data = 4'h4; //> 
    18'h15286: Data = 4'h4; //> 
    18'h15287: Data = 4'h4; //> 
    18'h15288: Data = 4'h7; //] 
    18'h15289: Data = 4'h2; //+ 
    18'h15290: Data = 4'h5; //< 
    18'h15291: Data = 4'h5; //< 
    18'h15292: Data = 4'h5; //< 
    18'h15293: Data = 4'h6; //[ 
    18'h15294: Data = 4'h3; //- 
    18'h15295: Data = 4'h4; //> 
    18'h15296: Data = 4'h4; //> 
    18'h15297: Data = 4'h4; //> 
    18'h15298: Data = 4'h3; //- 
    18'h15299: Data = 4'h4; //> 
    18'h15300: Data = 4'h6; //[ 
    18'h15301: Data = 4'h3; //- 
    18'h15302: Data = 4'h5; //< 
    18'h15303: Data = 4'h5; //< 
    18'h15304: Data = 4'h5; //< 
    18'h15305: Data = 4'h5; //< 
    18'h15306: Data = 4'h2; //+ 
    18'h15307: Data = 4'h4; //> 
    18'h15308: Data = 4'h4; //> 
    18'h15309: Data = 4'h4; //> 
    18'h15310: Data = 4'h4; //> 
    18'h15311: Data = 4'h7; //] 
    18'h15312: Data = 4'h5; //< 
    18'h15313: Data = 4'h5; //< 
    18'h15314: Data = 4'h5; //< 
    18'h15315: Data = 4'h5; //< 
    18'h15316: Data = 4'h6; //[ 
    18'h15317: Data = 4'h3; //- 
    18'h15318: Data = 4'h4; //> 
    18'h15319: Data = 4'h4; //> 
    18'h15320: Data = 4'h4; //> 
    18'h15321: Data = 4'h4; //> 
    18'h15322: Data = 4'h2; //+ 
    18'h15323: Data = 4'h5; //< 
    18'h15324: Data = 4'h5; //< 
    18'h15325: Data = 4'h5; //< 
    18'h15326: Data = 4'h5; //< 
    18'h15327: Data = 4'h5; //< 
    18'h15328: Data = 4'h5; //< 
    18'h15329: Data = 4'h5; //< 
    18'h15330: Data = 4'h5; //< 
    18'h15331: Data = 4'h5; //< 
    18'h15332: Data = 4'h5; //< 
    18'h15333: Data = 4'h5; //< 
    18'h15334: Data = 4'h5; //< 
    18'h15335: Data = 4'h5; //< 
    18'h15336: Data = 4'h6; //[ 
    18'h15337: Data = 4'h5; //< 
    18'h15338: Data = 4'h5; //< 
    18'h15339: Data = 4'h5; //< 
    18'h15340: Data = 4'h5; //< 
    18'h15341: Data = 4'h5; //< 
    18'h15342: Data = 4'h5; //< 
    18'h15343: Data = 4'h5; //< 
    18'h15344: Data = 4'h5; //< 
    18'h15345: Data = 4'h5; //< 
    18'h15346: Data = 4'h7; //] 
    18'h15347: Data = 4'h4; //> 
    18'h15348: Data = 4'h4; //> 
    18'h15349: Data = 4'h4; //> 
    18'h15350: Data = 4'h4; //> 
    18'h15351: Data = 4'ha; //0 
    18'h15352: Data = 4'h2; //+ 
    18'h15353: Data = 4'h4; //> 
    18'h15354: Data = 4'h4; //> 
    18'h15355: Data = 4'h4; //> 
    18'h15356: Data = 4'h4; //> 
    18'h15357: Data = 4'h4; //> 
    18'h15358: Data = 4'h6; //[ 
    18'h15359: Data = 4'h4; //> 
    18'h15360: Data = 4'h4; //> 
    18'h15361: Data = 4'h4; //> 
    18'h15362: Data = 4'h4; //> 
    18'h15363: Data = 4'h4; //> 
    18'h15364: Data = 4'h4; //> 
    18'h15365: Data = 4'h4; //> 
    18'h15366: Data = 4'h4; //> 
    18'h15367: Data = 4'h4; //> 
    18'h15368: Data = 4'h7; //] 
    18'h15369: Data = 4'h4; //> 
    18'h15370: Data = 4'h2; //+ 
    18'h15371: Data = 4'h5; //< 
    18'h15372: Data = 4'h7; //] 
    18'h15373: Data = 4'h7; //] 
    18'h15374: Data = 4'h2; //+ 
    18'h15375: Data = 4'h4; //> 
    18'h15376: Data = 4'h4; //> 
    18'h15377: Data = 4'h4; //> 
    18'h15378: Data = 4'h4; //> 
    18'h15379: Data = 4'h6; //[ 
    18'h15380: Data = 4'h3; //- 
    18'h15381: Data = 4'h5; //< 
    18'h15382: Data = 4'h5; //< 
    18'h15383: Data = 4'h5; //< 
    18'h15384: Data = 4'h5; //< 
    18'h15385: Data = 4'h3; //- 
    18'h15386: Data = 4'h4; //> 
    18'h15387: Data = 4'h4; //> 
    18'h15388: Data = 4'h4; //> 
    18'h15389: Data = 4'h4; //> 
    18'h15390: Data = 4'h7; //] 
    18'h15391: Data = 4'h2; //+ 
    18'h15392: Data = 4'h5; //< 
    18'h15393: Data = 4'h5; //< 
    18'h15394: Data = 4'h5; //< 
    18'h15395: Data = 4'h5; //< 
    18'h15396: Data = 4'h6; //[ 
    18'h15397: Data = 4'h3; //- 
    18'h15398: Data = 4'h4; //> 
    18'h15399: Data = 4'h4; //> 
    18'h15400: Data = 4'h4; //> 
    18'h15401: Data = 4'h4; //> 
    18'h15402: Data = 4'h3; //- 
    18'h15403: Data = 4'h5; //< 
    18'h15404: Data = 4'h6; //[ 
    18'h15405: Data = 4'h3; //- 
    18'h15406: Data = 4'h5; //< 
    18'h15407: Data = 4'h5; //< 
    18'h15408: Data = 4'h5; //< 
    18'h15409: Data = 4'h2; //+ 
    18'h15410: Data = 4'h4; //> 
    18'h15411: Data = 4'h4; //> 
    18'h15412: Data = 4'h4; //> 
    18'h15413: Data = 4'h7; //] 
    18'h15414: Data = 4'h5; //< 
    18'h15415: Data = 4'h5; //< 
    18'h15416: Data = 4'h5; //< 
    18'h15417: Data = 4'h6; //[ 
    18'h15418: Data = 4'h3; //- 
    18'h15419: Data = 4'h4; //> 
    18'h15420: Data = 4'h4; //> 
    18'h15421: Data = 4'h4; //> 
    18'h15422: Data = 4'h2; //+ 
    18'h15423: Data = 4'h5; //< 
    18'h15424: Data = 4'h5; //< 
    18'h15425: Data = 4'h5; //< 
    18'h15426: Data = 4'h5; //< 
    18'h15427: Data = 4'h5; //< 
    18'h15428: Data = 4'h5; //< 
    18'h15429: Data = 4'h5; //< 
    18'h15430: Data = 4'h5; //< 
    18'h15431: Data = 4'h5; //< 
    18'h15432: Data = 4'h5; //< 
    18'h15433: Data = 4'h5; //< 
    18'h15434: Data = 4'h5; //< 
    18'h15435: Data = 4'h6; //[ 
    18'h15436: Data = 4'h5; //< 
    18'h15437: Data = 4'h5; //< 
    18'h15438: Data = 4'h5; //< 
    18'h15439: Data = 4'h5; //< 
    18'h15440: Data = 4'h5; //< 
    18'h15441: Data = 4'h5; //< 
    18'h15442: Data = 4'h5; //< 
    18'h15443: Data = 4'h5; //< 
    18'h15444: Data = 4'h5; //< 
    18'h15445: Data = 4'h7; //] 
    18'h15446: Data = 4'h4; //> 
    18'h15447: Data = 4'h4; //> 
    18'h15448: Data = 4'h4; //> 
    18'h15449: Data = 4'ha; //0 
    18'h15450: Data = 4'h2; //+ 
    18'h15451: Data = 4'h4; //> 
    18'h15452: Data = 4'h4; //> 
    18'h15453: Data = 4'h4; //> 
    18'h15454: Data = 4'h4; //> 
    18'h15455: Data = 4'h4; //> 
    18'h15456: Data = 4'h4; //> 
    18'h15457: Data = 4'h6; //[ 
    18'h15458: Data = 4'h4; //> 
    18'h15459: Data = 4'h4; //> 
    18'h15460: Data = 4'h4; //> 
    18'h15461: Data = 4'h4; //> 
    18'h15462: Data = 4'h4; //> 
    18'h15463: Data = 4'h4; //> 
    18'h15464: Data = 4'h4; //> 
    18'h15465: Data = 4'h4; //> 
    18'h15466: Data = 4'h4; //> 
    18'h15467: Data = 4'h7; //] 
    18'h15468: Data = 4'h4; //> 
    18'h15469: Data = 4'ha; //0 
    18'h15470: Data = 4'h2; //+ 
    18'h15471: Data = 4'h5; //< 
    18'h15472: Data = 4'h7; //] 
    18'h15473: Data = 4'h7; //] 
    18'h15474: Data = 4'h2; //+ 
    18'h15475: Data = 4'h4; //> 
    18'h15476: Data = 4'h6; //[ 
    18'h15477: Data = 4'h3; //- 
    18'h15478: Data = 4'h5; //< 
    18'h15479: Data = 4'h6; //[ 
    18'h15480: Data = 4'h4; //> 
    18'h15481: Data = 4'h4; //> 
    18'h15482: Data = 4'h4; //> 
    18'h15483: Data = 4'h4; //> 
    18'h15484: Data = 4'h4; //> 
    18'h15485: Data = 4'h4; //> 
    18'h15486: Data = 4'h4; //> 
    18'h15487: Data = 4'h4; //> 
    18'h15488: Data = 4'h4; //> 
    18'h15489: Data = 4'h7; //] 
    18'h15490: Data = 4'h5; //< 
    18'h15491: Data = 4'h5; //< 
    18'h15492: Data = 4'h5; //< 
    18'h15493: Data = 4'h5; //< 
    18'h15494: Data = 4'h5; //< 
    18'h15495: Data = 4'h5; //< 
    18'h15496: Data = 4'h5; //< 
    18'h15497: Data = 4'h5; //< 
    18'h15498: Data = 4'h7; //] 
    18'h15499: Data = 4'h4; //> 
    18'h15500: Data = 4'h4; //> 
    18'h15501: Data = 4'h4; //> 
    18'h15502: Data = 4'h4; //> 
    18'h15503: Data = 4'h4; //> 
    18'h15504: Data = 4'h4; //> 
    18'h15505: Data = 4'h4; //> 
    18'h15506: Data = 4'h4; //> 
    18'h15507: Data = 4'h7; //] 
    18'h15508: Data = 4'h5; //< 
    18'h15509: Data = 4'h5; //< 
    18'h15510: Data = 4'h5; //< 
    18'h15511: Data = 4'h5; //< 
    18'h15512: Data = 4'h5; //< 
    18'h15513: Data = 4'h5; //< 
    18'h15514: Data = 4'h5; //< 
    18'h15515: Data = 4'h5; //< 
    18'h15516: Data = 4'h5; //< 
    18'h15517: Data = 4'h6; //[ 
    18'h15518: Data = 4'h5; //< 
    18'h15519: Data = 4'h5; //< 
    18'h15520: Data = 4'h5; //< 
    18'h15521: Data = 4'h5; //< 
    18'h15522: Data = 4'h5; //< 
    18'h15523: Data = 4'h5; //< 
    18'h15524: Data = 4'h5; //< 
    18'h15525: Data = 4'h5; //< 
    18'h15526: Data = 4'h5; //< 
    18'h15527: Data = 4'h7; //] 
    18'h15528: Data = 4'h4; //> 
    18'h15529: Data = 4'h4; //> 
    18'h15530: Data = 4'h4; //> 
    18'h15531: Data = 4'h6; //[ 
    18'h15532: Data = 4'h3; //- 
    18'h15533: Data = 4'h5; //< 
    18'h15534: Data = 4'h5; //< 
    18'h15535: Data = 4'h5; //< 
    18'h15536: Data = 4'h2; //+ 
    18'h15537: Data = 4'h4; //> 
    18'h15538: Data = 4'h4; //> 
    18'h15539: Data = 4'h4; //> 
    18'h15540: Data = 4'h7; //] 
    18'h15541: Data = 4'h5; //< 
    18'h15542: Data = 4'h5; //< 
    18'h15543: Data = 4'h5; //< 
    18'h15544: Data = 4'h6; //[ 
    18'h15545: Data = 4'h3; //- 
    18'h15546: Data = 4'h4; //> 
    18'h15547: Data = 4'h4; //> 
    18'h15548: Data = 4'h4; //> 
    18'h15549: Data = 4'h2; //+ 
    18'h15550: Data = 4'h4; //> 
    18'h15551: Data = 4'h4; //> 
    18'h15552: Data = 4'h4; //> 
    18'h15553: Data = 4'h4; //> 
    18'h15554: Data = 4'h4; //> 
    18'h15555: Data = 4'h4; //> 
    18'h15556: Data = 4'h6; //[ 
    18'h15557: Data = 4'h4; //> 
    18'h15558: Data = 4'h2; //+ 
    18'h15559: Data = 4'h4; //> 
    18'h15560: Data = 4'h4; //> 
    18'h15561: Data = 4'h4; //> 
    18'h15562: Data = 4'h6; //[ 
    18'h15563: Data = 4'h3; //- 
    18'h15564: Data = 4'h5; //< 
    18'h15565: Data = 4'h5; //< 
    18'h15566: Data = 4'h5; //< 
    18'h15567: Data = 4'h3; //- 
    18'h15568: Data = 4'h4; //> 
    18'h15569: Data = 4'h4; //> 
    18'h15570: Data = 4'h4; //> 
    18'h15571: Data = 4'h7; //] 
    18'h15572: Data = 4'h5; //< 
    18'h15573: Data = 4'h5; //< 
    18'h15574: Data = 4'h5; //< 
    18'h15575: Data = 4'h6; //[ 
    18'h15576: Data = 4'h3; //- 
    18'h15577: Data = 4'h4; //> 
    18'h15578: Data = 4'h4; //> 
    18'h15579: Data = 4'h4; //> 
    18'h15580: Data = 4'h2; //+ 
    18'h15581: Data = 4'h5; //< 
    18'h15582: Data = 4'h5; //< 
    18'h15583: Data = 4'h5; //< 
    18'h15584: Data = 4'h7; //] 
    18'h15585: Data = 4'h4; //> 
    18'h15586: Data = 4'h4; //> 
    18'h15587: Data = 4'h4; //> 
    18'h15588: Data = 4'h4; //> 
    18'h15589: Data = 4'h4; //> 
    18'h15590: Data = 4'h4; //> 
    18'h15591: Data = 4'h4; //> 
    18'h15592: Data = 4'h4; //> 
    18'h15593: Data = 4'h7; //] 
    18'h15594: Data = 4'h5; //< 
    18'h15595: Data = 4'h5; //< 
    18'h15596: Data = 4'h5; //< 
    18'h15597: Data = 4'h5; //< 
    18'h15598: Data = 4'h5; //< 
    18'h15599: Data = 4'h5; //< 
    18'h15600: Data = 4'h5; //< 
    18'h15601: Data = 4'h5; //< 
    18'h15602: Data = 4'h2; //+ 
    18'h15603: Data = 4'h5; //< 
    18'h15604: Data = 4'h6; //[ 
    18'h15605: Data = 4'h4; //> 
    18'h15606: Data = 4'h6; //[ 
    18'h15607: Data = 4'h3; //- 
    18'h15608: Data = 4'h4; //> 
    18'h15609: Data = 4'h2; //+ 
    18'h15610: Data = 4'h4; //> 
    18'h15611: Data = 4'h6; //[ 
    18'h15612: Data = 4'h3; //- 
    18'h15613: Data = 4'h5; //< 
    18'h15614: Data = 4'h3; //- 
    18'h15615: Data = 4'h5; //< 
    18'h15616: Data = 4'h5; //< 
    18'h15617: Data = 4'h5; //< 
    18'h15618: Data = 4'h5; //< 
    18'h15619: Data = 4'h5; //< 
    18'h15620: Data = 4'h5; //< 
    18'h15621: Data = 4'h5; //< 
    18'h15622: Data = 4'h5; //< 
    18'h15623: Data = 4'h5; //< 
    18'h15624: Data = 4'h5; //< 
    18'h15625: Data = 4'h2; //+ 
    18'h15626: Data = 4'h4; //> 
    18'h15627: Data = 4'h4; //> 
    18'h15628: Data = 4'h4; //> 
    18'h15629: Data = 4'h4; //> 
    18'h15630: Data = 4'h4; //> 
    18'h15631: Data = 4'h4; //> 
    18'h15632: Data = 4'h4; //> 
    18'h15633: Data = 4'h4; //> 
    18'h15634: Data = 4'h4; //> 
    18'h15635: Data = 4'h4; //> 
    18'h15636: Data = 4'h4; //> 
    18'h15637: Data = 4'h4; //> 
    18'h15638: Data = 4'h6; //[ 
    18'h15639: Data = 4'h3; //- 
    18'h15640: Data = 4'h5; //< 
    18'h15641: Data = 4'h5; //< 
    18'h15642: Data = 4'h2; //+ 
    18'h15643: Data = 4'h4; //> 
    18'h15644: Data = 4'h4; //> 
    18'h15645: Data = 4'h7; //] 
    18'h15646: Data = 4'h5; //< 
    18'h15647: Data = 4'h7; //] 
    18'h15648: Data = 4'h4; //> 
    18'h15649: Data = 4'h6; //[ 
    18'h15650: Data = 4'h3; //- 
    18'h15651: Data = 4'h5; //< 
    18'h15652: Data = 4'h5; //< 
    18'h15653: Data = 4'h3; //- 
    18'h15654: Data = 4'h5; //< 
    18'h15655: Data = 4'h5; //< 
    18'h15656: Data = 4'h5; //< 
    18'h15657: Data = 4'h5; //< 
    18'h15658: Data = 4'h5; //< 
    18'h15659: Data = 4'h5; //< 
    18'h15660: Data = 4'h5; //< 
    18'h15661: Data = 4'h5; //< 
    18'h15662: Data = 4'h5; //< 
    18'h15663: Data = 4'h5; //< 
    18'h15664: Data = 4'h2; //+ 
    18'h15665: Data = 4'h4; //> 
    18'h15666: Data = 4'h4; //> 
    18'h15667: Data = 4'h4; //> 
    18'h15668: Data = 4'h4; //> 
    18'h15669: Data = 4'h4; //> 
    18'h15670: Data = 4'h4; //> 
    18'h15671: Data = 4'h4; //> 
    18'h15672: Data = 4'h4; //> 
    18'h15673: Data = 4'h4; //> 
    18'h15674: Data = 4'h4; //> 
    18'h15675: Data = 4'h4; //> 
    18'h15676: Data = 4'h4; //> 
    18'h15677: Data = 4'h7; //] 
    18'h15678: Data = 4'h5; //< 
    18'h15679: Data = 4'h5; //< 
    18'h15680: Data = 4'h5; //< 
    18'h15681: Data = 4'h7; //] 
    18'h15682: Data = 4'h4; //> 
    18'h15683: Data = 4'h4; //> 
    18'h15684: Data = 4'h6; //[ 
    18'h15685: Data = 4'h3; //- 
    18'h15686: Data = 4'h5; //< 
    18'h15687: Data = 4'h2; //+ 
    18'h15688: Data = 4'h4; //> 
    18'h15689: Data = 4'h4; //> 
    18'h15690: Data = 4'h6; //[ 
    18'h15691: Data = 4'h3; //- 
    18'h15692: Data = 4'h5; //< 
    18'h15693: Data = 4'h5; //< 
    18'h15694: Data = 4'h3; //- 
    18'h15695: Data = 4'h5; //< 
    18'h15696: Data = 4'h5; //< 
    18'h15697: Data = 4'h5; //< 
    18'h15698: Data = 4'h5; //< 
    18'h15699: Data = 4'h5; //< 
    18'h15700: Data = 4'h5; //< 
    18'h15701: Data = 4'h5; //< 
    18'h15702: Data = 4'h5; //< 
    18'h15703: Data = 4'h5; //< 
    18'h15704: Data = 4'h5; //< 
    18'h15705: Data = 4'h2; //+ 
    18'h15706: Data = 4'h4; //> 
    18'h15707: Data = 4'h4; //> 
    18'h15708: Data = 4'h4; //> 
    18'h15709: Data = 4'h4; //> 
    18'h15710: Data = 4'h4; //> 
    18'h15711: Data = 4'h4; //> 
    18'h15712: Data = 4'h4; //> 
    18'h15713: Data = 4'h4; //> 
    18'h15714: Data = 4'h4; //> 
    18'h15715: Data = 4'h4; //> 
    18'h15716: Data = 4'h4; //> 
    18'h15717: Data = 4'h4; //> 
    18'h15718: Data = 4'h7; //] 
    18'h15719: Data = 4'h5; //< 
    18'h15720: Data = 4'h7; //] 
    18'h15721: Data = 4'h4; //> 
    18'h15722: Data = 4'h6; //[ 
    18'h15723: Data = 4'h3; //- 
    18'h15724: Data = 4'h5; //< 
    18'h15725: Data = 4'h5; //< 
    18'h15726: Data = 4'h2; //+ 
    18'h15727: Data = 4'h4; //> 
    18'h15728: Data = 4'h4; //> 
    18'h15729: Data = 4'h7; //] 
    18'h15730: Data = 4'h5; //< 
    18'h15731: Data = 4'h5; //< 
    18'h15732: Data = 4'h5; //< 
    18'h15733: Data = 4'h5; //< 
    18'h15734: Data = 4'h5; //< 
    18'h15735: Data = 4'h5; //< 
    18'h15736: Data = 4'h5; //< 
    18'h15737: Data = 4'h5; //< 
    18'h15738: Data = 4'h5; //< 
    18'h15739: Data = 4'h5; //< 
    18'h15740: Data = 4'h5; //< 
    18'h15741: Data = 4'h5; //< 
    18'h15742: Data = 4'h5; //< 
    18'h15743: Data = 4'h7; //] 
    18'h15744: Data = 4'h7; //] 
    18'h15745: Data = 4'h4; //> 
    18'h15746: Data = 4'h4; //> 
    18'h15747: Data = 4'h4; //> 
    18'h15748: Data = 4'h4; //> 
    18'h15749: Data = 4'h6; //[ 
    18'h15750: Data = 4'h3; //- 
    18'h15751: Data = 4'h5; //< 
    18'h15752: Data = 4'h5; //< 
    18'h15753: Data = 4'h5; //< 
    18'h15754: Data = 4'h5; //< 
    18'h15755: Data = 4'h2; //+ 
    18'h15756: Data = 4'h4; //> 
    18'h15757: Data = 4'h4; //> 
    18'h15758: Data = 4'h4; //> 
    18'h15759: Data = 4'h4; //> 
    18'h15760: Data = 4'h7; //] 
    18'h15761: Data = 4'h5; //< 
    18'h15762: Data = 4'h5; //< 
    18'h15763: Data = 4'h5; //< 
    18'h15764: Data = 4'h5; //< 
    18'h15765: Data = 4'h6; //[ 
    18'h15766: Data = 4'h3; //- 
    18'h15767: Data = 4'h4; //> 
    18'h15768: Data = 4'h4; //> 
    18'h15769: Data = 4'h4; //> 
    18'h15770: Data = 4'h4; //> 
    18'h15771: Data = 4'h2; //+ 
    18'h15772: Data = 4'h4; //> 
    18'h15773: Data = 4'h4; //> 
    18'h15774: Data = 4'h4; //> 
    18'h15775: Data = 4'h4; //> 
    18'h15776: Data = 4'h4; //> 
    18'h15777: Data = 4'h6; //[ 
    18'h15778: Data = 4'h4; //> 
    18'h15779: Data = 4'h2; //+ 
    18'h15780: Data = 4'h4; //> 
    18'h15781: Data = 4'h4; //> 
    18'h15782: Data = 4'h6; //[ 
    18'h15783: Data = 4'h3; //- 
    18'h15784: Data = 4'h5; //< 
    18'h15785: Data = 4'h5; //< 
    18'h15786: Data = 4'h3; //- 
    18'h15787: Data = 4'h4; //> 
    18'h15788: Data = 4'h4; //> 
    18'h15789: Data = 4'h7; //] 
    18'h15790: Data = 4'h5; //< 
    18'h15791: Data = 4'h5; //< 
    18'h15792: Data = 4'h6; //[ 
    18'h15793: Data = 4'h3; //- 
    18'h15794: Data = 4'h4; //> 
    18'h15795: Data = 4'h4; //> 
    18'h15796: Data = 4'h2; //+ 
    18'h15797: Data = 4'h5; //< 
    18'h15798: Data = 4'h5; //< 
    18'h15799: Data = 4'h7; //] 
    18'h15800: Data = 4'h4; //> 
    18'h15801: Data = 4'h4; //> 
    18'h15802: Data = 4'h4; //> 
    18'h15803: Data = 4'h4; //> 
    18'h15804: Data = 4'h4; //> 
    18'h15805: Data = 4'h4; //> 
    18'h15806: Data = 4'h4; //> 
    18'h15807: Data = 4'h4; //> 
    18'h15808: Data = 4'h7; //] 
    18'h15809: Data = 4'h5; //< 
    18'h15810: Data = 4'h5; //< 
    18'h15811: Data = 4'h5; //< 
    18'h15812: Data = 4'h5; //< 
    18'h15813: Data = 4'h5; //< 
    18'h15814: Data = 4'h5; //< 
    18'h15815: Data = 4'h5; //< 
    18'h15816: Data = 4'h5; //< 
    18'h15817: Data = 4'h2; //+ 
    18'h15818: Data = 4'h5; //< 
    18'h15819: Data = 4'h6; //[ 
    18'h15820: Data = 4'h4; //> 
    18'h15821: Data = 4'h6; //[ 
    18'h15822: Data = 4'h3; //- 
    18'h15823: Data = 4'h4; //> 
    18'h15824: Data = 4'h2; //+ 
    18'h15825: Data = 4'h4; //> 
    18'h15826: Data = 4'h4; //> 
    18'h15827: Data = 4'h6; //[ 
    18'h15828: Data = 4'h3; //- 
    18'h15829: Data = 4'h5; //< 
    18'h15830: Data = 4'h5; //< 
    18'h15831: Data = 4'h3; //- 
    18'h15832: Data = 4'h5; //< 
    18'h15833: Data = 4'h5; //< 
    18'h15834: Data = 4'h5; //< 
    18'h15835: Data = 4'h5; //< 
    18'h15836: Data = 4'h5; //< 
    18'h15837: Data = 4'h5; //< 
    18'h15838: Data = 4'h5; //< 
    18'h15839: Data = 4'h5; //< 
    18'h15840: Data = 4'h5; //< 
    18'h15841: Data = 4'h5; //< 
    18'h15842: Data = 4'h2; //+ 
    18'h15843: Data = 4'h4; //> 
    18'h15844: Data = 4'h4; //> 
    18'h15845: Data = 4'h4; //> 
    18'h15846: Data = 4'h4; //> 
    18'h15847: Data = 4'h4; //> 
    18'h15848: Data = 4'h4; //> 
    18'h15849: Data = 4'h4; //> 
    18'h15850: Data = 4'h4; //> 
    18'h15851: Data = 4'h4; //> 
    18'h15852: Data = 4'h4; //> 
    18'h15853: Data = 4'h4; //> 
    18'h15854: Data = 4'h6; //[ 
    18'h15855: Data = 4'h3; //- 
    18'h15856: Data = 4'h5; //< 
    18'h15857: Data = 4'h2; //+ 
    18'h15858: Data = 4'h4; //> 
    18'h15859: Data = 4'h7; //] 
    18'h15860: Data = 4'h4; //> 
    18'h15861: Data = 4'h7; //] 
    18'h15862: Data = 4'h5; //< 
    18'h15863: Data = 4'h6; //[ 
    18'h15864: Data = 4'h3; //- 
    18'h15865: Data = 4'h5; //< 
    18'h15866: Data = 4'h3; //- 
    18'h15867: Data = 4'h5; //< 
    18'h15868: Data = 4'h5; //< 
    18'h15869: Data = 4'h5; //< 
    18'h15870: Data = 4'h5; //< 
    18'h15871: Data = 4'h5; //< 
    18'h15872: Data = 4'h5; //< 
    18'h15873: Data = 4'h5; //< 
    18'h15874: Data = 4'h5; //< 
    18'h15875: Data = 4'h5; //< 
    18'h15876: Data = 4'h5; //< 
    18'h15877: Data = 4'h2; //+ 
    18'h15878: Data = 4'h4; //> 
    18'h15879: Data = 4'h4; //> 
    18'h15880: Data = 4'h4; //> 
    18'h15881: Data = 4'h4; //> 
    18'h15882: Data = 4'h4; //> 
    18'h15883: Data = 4'h4; //> 
    18'h15884: Data = 4'h4; //> 
    18'h15885: Data = 4'h4; //> 
    18'h15886: Data = 4'h4; //> 
    18'h15887: Data = 4'h4; //> 
    18'h15888: Data = 4'h4; //> 
    18'h15889: Data = 4'h7; //] 
    18'h15890: Data = 4'h5; //< 
    18'h15891: Data = 4'h5; //< 
    18'h15892: Data = 4'h7; //] 
    18'h15893: Data = 4'h4; //> 
    18'h15894: Data = 4'h4; //> 
    18'h15895: Data = 4'h4; //> 
    18'h15896: Data = 4'h6; //[ 
    18'h15897: Data = 4'h3; //- 
    18'h15898: Data = 4'h5; //< 
    18'h15899: Data = 4'h5; //< 
    18'h15900: Data = 4'h2; //+ 
    18'h15901: Data = 4'h4; //> 
    18'h15902: Data = 4'h6; //[ 
    18'h15903: Data = 4'h3; //- 
    18'h15904: Data = 4'h5; //< 
    18'h15905: Data = 4'h3; //- 
    18'h15906: Data = 4'h5; //< 
    18'h15907: Data = 4'h5; //< 
    18'h15908: Data = 4'h5; //< 
    18'h15909: Data = 4'h5; //< 
    18'h15910: Data = 4'h5; //< 
    18'h15911: Data = 4'h5; //< 
    18'h15912: Data = 4'h5; //< 
    18'h15913: Data = 4'h5; //< 
    18'h15914: Data = 4'h5; //< 
    18'h15915: Data = 4'h5; //< 
    18'h15916: Data = 4'h2; //+ 
    18'h15917: Data = 4'h4; //> 
    18'h15918: Data = 4'h4; //> 
    18'h15919: Data = 4'h4; //> 
    18'h15920: Data = 4'h4; //> 
    18'h15921: Data = 4'h4; //> 
    18'h15922: Data = 4'h4; //> 
    18'h15923: Data = 4'h4; //> 
    18'h15924: Data = 4'h4; //> 
    18'h15925: Data = 4'h4; //> 
    18'h15926: Data = 4'h4; //> 
    18'h15927: Data = 4'h4; //> 
    18'h15928: Data = 4'h7; //] 
    18'h15929: Data = 4'h4; //> 
    18'h15930: Data = 4'h7; //] 
    18'h15931: Data = 4'h5; //< 
    18'h15932: Data = 4'h6; //[ 
    18'h15933: Data = 4'h3; //- 
    18'h15934: Data = 4'h5; //< 
    18'h15935: Data = 4'h2; //+ 
    18'h15936: Data = 4'h4; //> 
    18'h15937: Data = 4'h7; //] 
    18'h15938: Data = 4'h5; //< 
    18'h15939: Data = 4'h5; //< 
    18'h15940: Data = 4'h5; //< 
    18'h15941: Data = 4'h5; //< 
    18'h15942: Data = 4'h5; //< 
    18'h15943: Data = 4'h5; //< 
    18'h15944: Data = 4'h5; //< 
    18'h15945: Data = 4'h5; //< 
    18'h15946: Data = 4'h5; //< 
    18'h15947: Data = 4'h5; //< 
    18'h15948: Data = 4'h5; //< 
    18'h15949: Data = 4'h5; //< 
    18'h15950: Data = 4'h7; //] 
    18'h15951: Data = 4'h4; //> 
    18'h15952: Data = 4'h4; //> 
    18'h15953: Data = 4'h4; //> 
    18'h15954: Data = 4'h4; //> 
    18'h15955: Data = 4'h4; //> 
    18'h15956: Data = 4'h2; //+ 
    18'h15957: Data = 4'h5; //< 
    18'h15958: Data = 4'h5; //< 
    18'h15959: Data = 4'h5; //< 
    18'h15960: Data = 4'h5; //< 
    18'h15961: Data = 4'h5; //< 
    18'h15962: Data = 4'h7; //] 
    18'h15963: Data = 4'h4; //> 
    18'h15964: Data = 4'h4; //> 
    18'h15965: Data = 4'h4; //> 
    18'h15966: Data = 4'h4; //> 
    18'h15967: Data = 4'h4; //> 
    18'h15968: Data = 4'h4; //> 
    18'h15969: Data = 4'h4; //> 
    18'h15970: Data = 4'h4; //> 
    18'h15971: Data = 4'h4; //> 
    18'h15972: Data = 4'h6; //[ 
    18'h15973: Data = 4'h4; //> 
    18'h15974: Data = 4'h4; //> 
    18'h15975: Data = 4'h4; //> 
    18'h15976: Data = 4'ha; //0 
    18'h15977: Data = 4'h4; //> 
    18'h15978: Data = 4'ha; //0 
    18'h15979: Data = 4'h4; //> 
    18'h15980: Data = 4'ha; //0 
    18'h15981: Data = 4'h4; //> 
    18'h15982: Data = 4'h4; //> 
    18'h15983: Data = 4'h4; //> 
    18'h15984: Data = 4'h4; //> 
    18'h15985: Data = 4'h7; //] 
    18'h15986: Data = 4'h5; //< 
    18'h15987: Data = 4'h5; //< 
    18'h15988: Data = 4'h5; //< 
    18'h15989: Data = 4'h5; //< 
    18'h15990: Data = 4'h5; //< 
    18'h15991: Data = 4'h5; //< 
    18'h15992: Data = 4'h5; //< 
    18'h15993: Data = 4'h5; //< 
    18'h15994: Data = 4'h5; //< 
    18'h15995: Data = 4'h6; //[ 
    18'h15996: Data = 4'h5; //< 
    18'h15997: Data = 4'h5; //< 
    18'h15998: Data = 4'h5; //< 
    18'h15999: Data = 4'h5; //< 
    18'h16000: Data = 4'h5; //< 
    18'h16001: Data = 4'h5; //< 
    18'h16002: Data = 4'h5; //< 
    18'h16003: Data = 4'h5; //< 
    18'h16004: Data = 4'h5; //< 
    18'h16005: Data = 4'h7; //] 
    18'h16006: Data = 4'h4; //> 
    18'h16007: Data = 4'h4; //> 
    18'h16008: Data = 4'h4; //> 
    18'h16009: Data = 4'ha; //0 
    18'h16010: Data = 4'h4; //> 
    18'h16011: Data = 4'ha; //0 
    18'h16012: Data = 4'h4; //> 
    18'h16013: Data = 4'h4; //> 
    18'h16014: Data = 4'h4; //> 
    18'h16015: Data = 4'h4; //> 
    18'h16016: Data = 4'h4; //> 
    18'h16017: Data = 4'h6; //[ 
    18'h16018: Data = 4'h4; //> 
    18'h16019: Data = 4'h4; //> 
    18'h16020: Data = 4'h4; //> 
    18'h16021: Data = 4'h4; //> 
    18'h16022: Data = 4'h4; //> 
    18'h16023: Data = 4'h4; //> 
    18'h16024: Data = 4'h4; //> 
    18'h16025: Data = 4'h6; //[ 
    18'h16026: Data = 4'h3; //- 
    18'h16027: Data = 4'h5; //< 
    18'h16028: Data = 4'h5; //< 
    18'h16029: Data = 4'h5; //< 
    18'h16030: Data = 4'h5; //< 
    18'h16031: Data = 4'h5; //< 
    18'h16032: Data = 4'h5; //< 
    18'h16033: Data = 4'h2; //+ 
    18'h16034: Data = 4'h4; //> 
    18'h16035: Data = 4'h4; //> 
    18'h16036: Data = 4'h4; //> 
    18'h16037: Data = 4'h4; //> 
    18'h16038: Data = 4'h4; //> 
    18'h16039: Data = 4'h4; //> 
    18'h16040: Data = 4'h7; //] 
    18'h16041: Data = 4'h5; //< 
    18'h16042: Data = 4'h5; //< 
    18'h16043: Data = 4'h5; //< 
    18'h16044: Data = 4'h5; //< 
    18'h16045: Data = 4'h5; //< 
    18'h16046: Data = 4'h5; //< 
    18'h16047: Data = 4'h6; //[ 
    18'h16048: Data = 4'h3; //- 
    18'h16049: Data = 4'h4; //> 
    18'h16050: Data = 4'h4; //> 
    18'h16051: Data = 4'h4; //> 
    18'h16052: Data = 4'h4; //> 
    18'h16053: Data = 4'h4; //> 
    18'h16054: Data = 4'h4; //> 
    18'h16055: Data = 4'h2; //+ 
    18'h16056: Data = 4'h5; //< 
    18'h16057: Data = 4'h5; //< 
    18'h16058: Data = 4'h5; //< 
    18'h16059: Data = 4'h5; //< 
    18'h16060: Data = 4'h2; //+ 
    18'h16061: Data = 4'h5; //< 
    18'h16062: Data = 4'h5; //< 
    18'h16063: Data = 4'h7; //] 
    18'h16064: Data = 4'h4; //> 
    18'h16065: Data = 4'h4; //> 
    18'h16066: Data = 4'h4; //> 
    18'h16067: Data = 4'h4; //> 
    18'h16068: Data = 4'h4; //> 
    18'h16069: Data = 4'h4; //> 
    18'h16070: Data = 4'h4; //> 
    18'h16071: Data = 4'h4; //> 
    18'h16072: Data = 4'h7; //] 
    18'h16073: Data = 4'h5; //< 
    18'h16074: Data = 4'h5; //< 
    18'h16075: Data = 4'h5; //< 
    18'h16076: Data = 4'h5; //< 
    18'h16077: Data = 4'h5; //< 
    18'h16078: Data = 4'h5; //< 
    18'h16079: Data = 4'h5; //< 
    18'h16080: Data = 4'h5; //< 
    18'h16081: Data = 4'h5; //< 
    18'h16082: Data = 4'h6; //[ 
    18'h16083: Data = 4'h5; //< 
    18'h16084: Data = 4'h5; //< 
    18'h16085: Data = 4'h5; //< 
    18'h16086: Data = 4'h5; //< 
    18'h16087: Data = 4'h5; //< 
    18'h16088: Data = 4'h5; //< 
    18'h16089: Data = 4'h5; //< 
    18'h16090: Data = 4'h5; //< 
    18'h16091: Data = 4'h5; //< 
    18'h16092: Data = 4'h7; //] 
    18'h16093: Data = 4'h4; //> 
    18'h16094: Data = 4'h4; //> 
    18'h16095: Data = 4'h4; //> 
    18'h16096: Data = 4'h4; //> 
    18'h16097: Data = 4'h2; //+ 
    18'h16098: Data = 4'h4; //> 
    18'h16099: Data = 4'h6; //[ 
    18'h16100: Data = 4'h3; //- 
    18'h16101: Data = 4'h5; //< 
    18'h16102: Data = 4'h3; //- 
    18'h16103: Data = 4'h5; //< 
    18'h16104: Data = 4'h5; //< 
    18'h16105: Data = 4'h5; //< 
    18'h16106: Data = 4'h5; //< 
    18'h16107: Data = 4'h2; //+ 
    18'h16108: Data = 4'h4; //> 
    18'h16109: Data = 4'h4; //> 
    18'h16110: Data = 4'h4; //> 
    18'h16111: Data = 4'h4; //> 
    18'h16112: Data = 4'h4; //> 
    18'h16113: Data = 4'h7; //] 
    18'h16114: Data = 4'h4; //> 
    18'h16115: Data = 4'h4; //> 
    18'h16116: Data = 4'h6; //[ 
    18'h16117: Data = 4'h3; //- 
    18'h16118: Data = 4'h5; //< 
    18'h16119: Data = 4'h5; //< 
    18'h16120: Data = 4'h5; //< 
    18'h16121: Data = 4'h5; //< 
    18'h16122: Data = 4'h5; //< 
    18'h16123: Data = 4'h5; //< 
    18'h16124: Data = 4'h5; //< 
    18'h16125: Data = 4'h6; //[ 
    18'h16126: Data = 4'h3; //- 
    18'h16127: Data = 4'h4; //> 
    18'h16128: Data = 4'h4; //> 
    18'h16129: Data = 4'h4; //> 
    18'h16130: Data = 4'h4; //> 
    18'h16131: Data = 4'h4; //> 
    18'h16132: Data = 4'h2; //+ 
    18'h16133: Data = 4'h5; //< 
    18'h16134: Data = 4'h2; //+ 
    18'h16135: Data = 4'h2; //+ 
    18'h16136: Data = 4'h5; //< 
    18'h16137: Data = 4'h5; //< 
    18'h16138: Data = 4'h5; //< 
    18'h16139: Data = 4'h5; //< 
    18'h16140: Data = 4'h7; //] 
    18'h16141: Data = 4'h4; //> 
    18'h16142: Data = 4'h4; //> 
    18'h16143: Data = 4'h4; //> 
    18'h16144: Data = 4'h4; //> 
    18'h16145: Data = 4'h4; //> 
    18'h16146: Data = 4'h6; //[ 
    18'h16147: Data = 4'h3; //- 
    18'h16148: Data = 4'h5; //< 
    18'h16149: Data = 4'h5; //< 
    18'h16150: Data = 4'h5; //< 
    18'h16151: Data = 4'h5; //< 
    18'h16152: Data = 4'h5; //< 
    18'h16153: Data = 4'h2; //+ 
    18'h16154: Data = 4'h4; //> 
    18'h16155: Data = 4'h4; //> 
    18'h16156: Data = 4'h4; //> 
    18'h16157: Data = 4'h4; //> 
    18'h16158: Data = 4'h4; //> 
    18'h16159: Data = 4'h7; //] 
    18'h16160: Data = 4'h5; //< 
    18'h16161: Data = 4'h3; //- 
    18'h16162: Data = 4'h4; //> 
    18'h16163: Data = 4'h2; //+ 
    18'h16164: Data = 4'h4; //> 
    18'h16165: Data = 4'h4; //> 
    18'h16166: Data = 4'h7; //] 
    18'h16167: Data = 4'h5; //< 
    18'h16168: Data = 4'h5; //< 
    18'h16169: Data = 4'h6; //[ 
    18'h16170: Data = 4'h3; //- 
    18'h16171: Data = 4'h4; //> 
    18'h16172: Data = 4'h4; //> 
    18'h16173: Data = 4'h2; //+ 
    18'h16174: Data = 4'h5; //< 
    18'h16175: Data = 4'h5; //< 
    18'h16176: Data = 4'h7; //] 
    18'h16177: Data = 4'h5; //< 
    18'h16178: Data = 4'h5; //< 
    18'h16179: Data = 4'h5; //< 
    18'h16180: Data = 4'h5; //< 
    18'h16181: Data = 4'h5; //< 
    18'h16182: Data = 4'h6; //[ 
    18'h16183: Data = 4'h3; //- 
    18'h16184: Data = 4'h4; //> 
    18'h16185: Data = 4'h4; //> 
    18'h16186: Data = 4'h4; //> 
    18'h16187: Data = 4'h4; //> 
    18'h16188: Data = 4'h4; //> 
    18'h16189: Data = 4'h2; //+ 
    18'h16190: Data = 4'h5; //< 
    18'h16191: Data = 4'h5; //< 
    18'h16192: Data = 4'h5; //< 
    18'h16193: Data = 4'h5; //< 
    18'h16194: Data = 4'h5; //< 
    18'h16195: Data = 4'h7; //] 
    18'h16196: Data = 4'h2; //+ 
    18'h16197: Data = 4'h4; //> 
    18'h16198: Data = 4'h4; //> 
    18'h16199: Data = 4'h4; //> 
    18'h16200: Data = 4'h4; //> 
    18'h16201: Data = 4'h6; //[ 
    18'h16202: Data = 4'h3; //- 
    18'h16203: Data = 4'h5; //< 
    18'h16204: Data = 4'h5; //< 
    18'h16205: Data = 4'h5; //< 
    18'h16206: Data = 4'h5; //< 
    18'h16207: Data = 4'h3; //- 
    18'h16208: Data = 4'h4; //> 
    18'h16209: Data = 4'h4; //> 
    18'h16210: Data = 4'h4; //> 
    18'h16211: Data = 4'h4; //> 
    18'h16212: Data = 4'h7; //] 
    18'h16213: Data = 4'h2; //+ 
    18'h16214: Data = 4'h5; //< 
    18'h16215: Data = 4'h5; //< 
    18'h16216: Data = 4'h5; //< 
    18'h16217: Data = 4'h5; //< 
    18'h16218: Data = 4'h6; //[ 
    18'h16219: Data = 4'h3; //- 
    18'h16220: Data = 4'h4; //> 
    18'h16221: Data = 4'h4; //> 
    18'h16222: Data = 4'h4; //> 
    18'h16223: Data = 4'h4; //> 
    18'h16224: Data = 4'h3; //- 
    18'h16225: Data = 4'h4; //> 
    18'h16226: Data = 4'h4; //> 
    18'h16227: Data = 4'h4; //> 
    18'h16228: Data = 4'h4; //> 
    18'h16229: Data = 4'h4; //> 
    18'h16230: Data = 4'h6; //[ 
    18'h16231: Data = 4'h4; //> 
    18'h16232: Data = 4'h4; //> 
    18'h16233: Data = 4'h4; //> 
    18'h16234: Data = 4'h6; //[ 
    18'h16235: Data = 4'h3; //- 
    18'h16236: Data = 4'h5; //< 
    18'h16237: Data = 4'h5; //< 
    18'h16238: Data = 4'h5; //< 
    18'h16239: Data = 4'h3; //- 
    18'h16240: Data = 4'h4; //> 
    18'h16241: Data = 4'h4; //> 
    18'h16242: Data = 4'h4; //> 
    18'h16243: Data = 4'h7; //] 
    18'h16244: Data = 4'h2; //+ 
    18'h16245: Data = 4'h5; //< 
    18'h16246: Data = 4'h5; //< 
    18'h16247: Data = 4'h5; //< 
    18'h16248: Data = 4'h6; //[ 
    18'h16249: Data = 4'h3; //- 
    18'h16250: Data = 4'h4; //> 
    18'h16251: Data = 4'h4; //> 
    18'h16252: Data = 4'h4; //> 
    18'h16253: Data = 4'h3; //- 
    18'h16254: Data = 4'h5; //< 
    18'h16255: Data = 4'h6; //[ 
    18'h16256: Data = 4'h3; //- 
    18'h16257: Data = 4'h5; //< 
    18'h16258: Data = 4'h5; //< 
    18'h16259: Data = 4'h2; //+ 
    18'h16260: Data = 4'h4; //> 
    18'h16261: Data = 4'h4; //> 
    18'h16262: Data = 4'h7; //] 
    18'h16263: Data = 4'h5; //< 
    18'h16264: Data = 4'h5; //< 
    18'h16265: Data = 4'h6; //[ 
    18'h16266: Data = 4'h3; //- 
    18'h16267: Data = 4'h4; //> 
    18'h16268: Data = 4'h4; //> 
    18'h16269: Data = 4'h2; //+ 
    18'h16270: Data = 4'h5; //< 
    18'h16271: Data = 4'h5; //< 
    18'h16272: Data = 4'h5; //< 
    18'h16273: Data = 4'h5; //< 
    18'h16274: Data = 4'h5; //< 
    18'h16275: Data = 4'h5; //< 
    18'h16276: Data = 4'h5; //< 
    18'h16277: Data = 4'h5; //< 
    18'h16278: Data = 4'h5; //< 
    18'h16279: Data = 4'h5; //< 
    18'h16280: Data = 4'h5; //< 
    18'h16281: Data = 4'h6; //[ 
    18'h16282: Data = 4'h5; //< 
    18'h16283: Data = 4'h5; //< 
    18'h16284: Data = 4'h5; //< 
    18'h16285: Data = 4'h5; //< 
    18'h16286: Data = 4'h5; //< 
    18'h16287: Data = 4'h5; //< 
    18'h16288: Data = 4'h5; //< 
    18'h16289: Data = 4'h5; //< 
    18'h16290: Data = 4'h5; //< 
    18'h16291: Data = 4'h7; //] 
    18'h16292: Data = 4'h4; //> 
    18'h16293: Data = 4'h4; //> 
    18'h16294: Data = 4'h4; //> 
    18'h16295: Data = 4'h4; //> 
    18'h16296: Data = 4'ha; //0 
    18'h16297: Data = 4'h2; //+ 
    18'h16298: Data = 4'h4; //> 
    18'h16299: Data = 4'h4; //> 
    18'h16300: Data = 4'h4; //> 
    18'h16301: Data = 4'h4; //> 
    18'h16302: Data = 4'h4; //> 
    18'h16303: Data = 4'h6; //[ 
    18'h16304: Data = 4'h4; //> 
    18'h16305: Data = 4'h4; //> 
    18'h16306: Data = 4'h4; //> 
    18'h16307: Data = 4'h4; //> 
    18'h16308: Data = 4'h4; //> 
    18'h16309: Data = 4'h4; //> 
    18'h16310: Data = 4'h4; //> 
    18'h16311: Data = 4'h4; //> 
    18'h16312: Data = 4'h4; //> 
    18'h16313: Data = 4'h7; //] 
    18'h16314: Data = 4'h4; //> 
    18'h16315: Data = 4'h2; //+ 
    18'h16316: Data = 4'h5; //< 
    18'h16317: Data = 4'h7; //] 
    18'h16318: Data = 4'h7; //] 
    18'h16319: Data = 4'h2; //+ 
    18'h16320: Data = 4'h4; //> 
    18'h16321: Data = 4'h4; //> 
    18'h16322: Data = 4'h6; //[ 
    18'h16323: Data = 4'h3; //- 
    18'h16324: Data = 4'h5; //< 
    18'h16325: Data = 4'h5; //< 
    18'h16326: Data = 4'h3; //- 
    18'h16327: Data = 4'h4; //> 
    18'h16328: Data = 4'h4; //> 
    18'h16329: Data = 4'h7; //] 
    18'h16330: Data = 4'h2; //+ 
    18'h16331: Data = 4'h5; //< 
    18'h16332: Data = 4'h5; //< 
    18'h16333: Data = 4'h6; //[ 
    18'h16334: Data = 4'h3; //- 
    18'h16335: Data = 4'h4; //> 
    18'h16336: Data = 4'h4; //> 
    18'h16337: Data = 4'h3; //- 
    18'h16338: Data = 4'h4; //> 
    18'h16339: Data = 4'h6; //[ 
    18'h16340: Data = 4'h3; //- 
    18'h16341: Data = 4'h5; //< 
    18'h16342: Data = 4'h5; //< 
    18'h16343: Data = 4'h5; //< 
    18'h16344: Data = 4'h2; //+ 
    18'h16345: Data = 4'h4; //> 
    18'h16346: Data = 4'h4; //> 
    18'h16347: Data = 4'h4; //> 
    18'h16348: Data = 4'h7; //] 
    18'h16349: Data = 4'h5; //< 
    18'h16350: Data = 4'h5; //< 
    18'h16351: Data = 4'h5; //< 
    18'h16352: Data = 4'h6; //[ 
    18'h16353: Data = 4'h3; //- 
    18'h16354: Data = 4'h4; //> 
    18'h16355: Data = 4'h4; //> 
    18'h16356: Data = 4'h4; //> 
    18'h16357: Data = 4'h2; //+ 
    18'h16358: Data = 4'h5; //< 
    18'h16359: Data = 4'h5; //< 
    18'h16360: Data = 4'h5; //< 
    18'h16361: Data = 4'h5; //< 
    18'h16362: Data = 4'h5; //< 
    18'h16363: Data = 4'h5; //< 
    18'h16364: Data = 4'h5; //< 
    18'h16365: Data = 4'h5; //< 
    18'h16366: Data = 4'h5; //< 
    18'h16367: Data = 4'h5; //< 
    18'h16368: Data = 4'h5; //< 
    18'h16369: Data = 4'h5; //< 
    18'h16370: Data = 4'h6; //[ 
    18'h16371: Data = 4'h5; //< 
    18'h16372: Data = 4'h5; //< 
    18'h16373: Data = 4'h5; //< 
    18'h16374: Data = 4'h5; //< 
    18'h16375: Data = 4'h5; //< 
    18'h16376: Data = 4'h5; //< 
    18'h16377: Data = 4'h5; //< 
    18'h16378: Data = 4'h5; //< 
    18'h16379: Data = 4'h5; //< 
    18'h16380: Data = 4'h7; //] 
    18'h16381: Data = 4'h4; //> 
    18'h16382: Data = 4'h4; //> 
    18'h16383: Data = 4'h4; //> 
    18'h16384: Data = 4'ha; //0 
    18'h16385: Data = 4'h2; //+ 
    18'h16386: Data = 4'h4; //> 
    18'h16387: Data = 4'h4; //> 
    18'h16388: Data = 4'h4; //> 
    18'h16389: Data = 4'h4; //> 
    18'h16390: Data = 4'h4; //> 
    18'h16391: Data = 4'h4; //> 
    18'h16392: Data = 4'h6; //[ 
    18'h16393: Data = 4'h4; //> 
    18'h16394: Data = 4'h4; //> 
    18'h16395: Data = 4'h4; //> 
    18'h16396: Data = 4'h4; //> 
    18'h16397: Data = 4'h4; //> 
    18'h16398: Data = 4'h4; //> 
    18'h16399: Data = 4'h4; //> 
    18'h16400: Data = 4'h4; //> 
    18'h16401: Data = 4'h4; //> 
    18'h16402: Data = 4'h7; //] 
    18'h16403: Data = 4'h4; //> 
    18'h16404: Data = 4'ha; //0 
    18'h16405: Data = 4'h2; //+ 
    18'h16406: Data = 4'h5; //< 
    18'h16407: Data = 4'h7; //] 
    18'h16408: Data = 4'h7; //] 
    18'h16409: Data = 4'h2; //+ 
    18'h16410: Data = 4'h4; //> 
    18'h16411: Data = 4'h6; //[ 
    18'h16412: Data = 4'h3; //- 
    18'h16413: Data = 4'h5; //< 
    18'h16414: Data = 4'h6; //[ 
    18'h16415: Data = 4'h4; //> 
    18'h16416: Data = 4'h4; //> 
    18'h16417: Data = 4'h4; //> 
    18'h16418: Data = 4'h4; //> 
    18'h16419: Data = 4'h4; //> 
    18'h16420: Data = 4'h4; //> 
    18'h16421: Data = 4'h4; //> 
    18'h16422: Data = 4'h4; //> 
    18'h16423: Data = 4'h4; //> 
    18'h16424: Data = 4'h7; //] 
    18'h16425: Data = 4'h5; //< 
    18'h16426: Data = 4'h5; //< 
    18'h16427: Data = 4'h5; //< 
    18'h16428: Data = 4'h5; //< 
    18'h16429: Data = 4'h5; //< 
    18'h16430: Data = 4'h5; //< 
    18'h16431: Data = 4'h5; //< 
    18'h16432: Data = 4'h5; //< 
    18'h16433: Data = 4'h7; //] 
    18'h16434: Data = 4'h4; //> 
    18'h16435: Data = 4'h4; //> 
    18'h16436: Data = 4'h4; //> 
    18'h16437: Data = 4'h4; //> 
    18'h16438: Data = 4'h4; //> 
    18'h16439: Data = 4'h4; //> 
    18'h16440: Data = 4'h4; //> 
    18'h16441: Data = 4'h4; //> 
    18'h16442: Data = 4'h7; //] 
    18'h16443: Data = 4'h5; //< 
    18'h16444: Data = 4'h5; //< 
    18'h16445: Data = 4'h5; //< 
    18'h16446: Data = 4'h5; //< 
    18'h16447: Data = 4'h5; //< 
    18'h16448: Data = 4'h5; //< 
    18'h16449: Data = 4'h5; //< 
    18'h16450: Data = 4'h5; //< 
    18'h16451: Data = 4'h5; //< 
    18'h16452: Data = 4'h6; //[ 
    18'h16453: Data = 4'h5; //< 
    18'h16454: Data = 4'h5; //< 
    18'h16455: Data = 4'h5; //< 
    18'h16456: Data = 4'h5; //< 
    18'h16457: Data = 4'h5; //< 
    18'h16458: Data = 4'h5; //< 
    18'h16459: Data = 4'h5; //< 
    18'h16460: Data = 4'h5; //< 
    18'h16461: Data = 4'h5; //< 
    18'h16462: Data = 4'h7; //] 
    18'h16463: Data = 4'h4; //> 
    18'h16464: Data = 4'h4; //> 
    18'h16465: Data = 4'h4; //> 
    18'h16466: Data = 4'h6; //[ 
    18'h16467: Data = 4'h3; //- 
    18'h16468: Data = 4'h5; //< 
    18'h16469: Data = 4'h5; //< 
    18'h16470: Data = 4'h5; //< 
    18'h16471: Data = 4'h2; //+ 
    18'h16472: Data = 4'h4; //> 
    18'h16473: Data = 4'h4; //> 
    18'h16474: Data = 4'h4; //> 
    18'h16475: Data = 4'h7; //] 
    18'h16476: Data = 4'h5; //< 
    18'h16477: Data = 4'h5; //< 
    18'h16478: Data = 4'h5; //< 
    18'h16479: Data = 4'h6; //[ 
    18'h16480: Data = 4'h3; //- 
    18'h16481: Data = 4'h4; //> 
    18'h16482: Data = 4'h4; //> 
    18'h16483: Data = 4'h4; //> 
    18'h16484: Data = 4'h2; //+ 
    18'h16485: Data = 4'h4; //> 
    18'h16486: Data = 4'h4; //> 
    18'h16487: Data = 4'h4; //> 
    18'h16488: Data = 4'h4; //> 
    18'h16489: Data = 4'h4; //> 
    18'h16490: Data = 4'h4; //> 
    18'h16491: Data = 4'h6; //[ 
    18'h16492: Data = 4'h4; //> 
    18'h16493: Data = 4'h2; //+ 
    18'h16494: Data = 4'h4; //> 
    18'h16495: Data = 4'h6; //[ 
    18'h16496: Data = 4'h3; //- 
    18'h16497: Data = 4'h5; //< 
    18'h16498: Data = 4'h3; //- 
    18'h16499: Data = 4'h4; //> 
    18'h16500: Data = 4'h7; //] 
    18'h16501: Data = 4'h5; //< 
    18'h16502: Data = 4'h6; //[ 
    18'h16503: Data = 4'h3; //- 
    18'h16504: Data = 4'h4; //> 
    18'h16505: Data = 4'h2; //+ 
    18'h16506: Data = 4'h5; //< 
    18'h16507: Data = 4'h7; //] 
    18'h16508: Data = 4'h4; //> 
    18'h16509: Data = 4'h4; //> 
    18'h16510: Data = 4'h4; //> 
    18'h16511: Data = 4'h4; //> 
    18'h16512: Data = 4'h4; //> 
    18'h16513: Data = 4'h4; //> 
    18'h16514: Data = 4'h4; //> 
    18'h16515: Data = 4'h4; //> 
    18'h16516: Data = 4'h7; //] 
    18'h16517: Data = 4'h5; //< 
    18'h16518: Data = 4'h5; //< 
    18'h16519: Data = 4'h5; //< 
    18'h16520: Data = 4'h5; //< 
    18'h16521: Data = 4'h5; //< 
    18'h16522: Data = 4'h5; //< 
    18'h16523: Data = 4'h5; //< 
    18'h16524: Data = 4'h5; //< 
    18'h16525: Data = 4'h2; //+ 
    18'h16526: Data = 4'h5; //< 
    18'h16527: Data = 4'h6; //[ 
    18'h16528: Data = 4'h4; //> 
    18'h16529: Data = 4'h6; //[ 
    18'h16530: Data = 4'h3; //- 
    18'h16531: Data = 4'h4; //> 
    18'h16532: Data = 4'h4; //> 
    18'h16533: Data = 4'h4; //> 
    18'h16534: Data = 4'h4; //> 
    18'h16535: Data = 4'h2; //+ 
    18'h16536: Data = 4'h5; //< 
    18'h16537: Data = 4'h5; //< 
    18'h16538: Data = 4'h6; //[ 
    18'h16539: Data = 4'h3; //- 
    18'h16540: Data = 4'h4; //> 
    18'h16541: Data = 4'h4; //> 
    18'h16542: Data = 4'h3; //- 
    18'h16543: Data = 4'h5; //< 
    18'h16544: Data = 4'h5; //< 
    18'h16545: Data = 4'h5; //< 
    18'h16546: Data = 4'h5; //< 
    18'h16547: Data = 4'h5; //< 
    18'h16548: Data = 4'h5; //< 
    18'h16549: Data = 4'h5; //< 
    18'h16550: Data = 4'h5; //< 
    18'h16551: Data = 4'h5; //< 
    18'h16552: Data = 4'h5; //< 
    18'h16553: Data = 4'h5; //< 
    18'h16554: Data = 4'h5; //< 
    18'h16555: Data = 4'h5; //< 
    18'h16556: Data = 4'h2; //+ 
    18'h16557: Data = 4'h4; //> 
    18'h16558: Data = 4'h4; //> 
    18'h16559: Data = 4'h4; //> 
    18'h16560: Data = 4'h4; //> 
    18'h16561: Data = 4'h4; //> 
    18'h16562: Data = 4'h4; //> 
    18'h16563: Data = 4'h4; //> 
    18'h16564: Data = 4'h4; //> 
    18'h16565: Data = 4'h4; //> 
    18'h16566: Data = 4'h4; //> 
    18'h16567: Data = 4'h6; //[ 
    18'h16568: Data = 4'h3; //- 
    18'h16569: Data = 4'h4; //> 
    18'h16570: Data = 4'h4; //> 
    18'h16571: Data = 4'h4; //> 
    18'h16572: Data = 4'h2; //+ 
    18'h16573: Data = 4'h5; //< 
    18'h16574: Data = 4'h5; //< 
    18'h16575: Data = 4'h5; //< 
    18'h16576: Data = 4'h7; //] 
    18'h16577: Data = 4'h4; //> 
    18'h16578: Data = 4'h7; //] 
    18'h16579: Data = 4'h5; //< 
    18'h16580: Data = 4'h6; //[ 
    18'h16581: Data = 4'h3; //- 
    18'h16582: Data = 4'h4; //> 
    18'h16583: Data = 4'h4; //> 
    18'h16584: Data = 4'h4; //> 
    18'h16585: Data = 4'h3; //- 
    18'h16586: Data = 4'h5; //< 
    18'h16587: Data = 4'h5; //< 
    18'h16588: Data = 4'h5; //< 
    18'h16589: Data = 4'h5; //< 
    18'h16590: Data = 4'h5; //< 
    18'h16591: Data = 4'h5; //< 
    18'h16592: Data = 4'h5; //< 
    18'h16593: Data = 4'h5; //< 
    18'h16594: Data = 4'h5; //< 
    18'h16595: Data = 4'h5; //< 
    18'h16596: Data = 4'h5; //< 
    18'h16597: Data = 4'h5; //< 
    18'h16598: Data = 4'h5; //< 
    18'h16599: Data = 4'h2; //+ 
    18'h16600: Data = 4'h4; //> 
    18'h16601: Data = 4'h4; //> 
    18'h16602: Data = 4'h4; //> 
    18'h16603: Data = 4'h4; //> 
    18'h16604: Data = 4'h4; //> 
    18'h16605: Data = 4'h4; //> 
    18'h16606: Data = 4'h4; //> 
    18'h16607: Data = 4'h4; //> 
    18'h16608: Data = 4'h4; //> 
    18'h16609: Data = 4'h4; //> 
    18'h16610: Data = 4'h7; //] 
    18'h16611: Data = 4'h5; //< 
    18'h16612: Data = 4'h7; //] 
    18'h16613: Data = 4'h4; //> 
    18'h16614: Data = 4'h4; //> 
    18'h16615: Data = 4'h6; //[ 
    18'h16616: Data = 4'h3; //- 
    18'h16617: Data = 4'h4; //> 
    18'h16618: Data = 4'h4; //> 
    18'h16619: Data = 4'h2; //+ 
    18'h16620: Data = 4'h5; //< 
    18'h16621: Data = 4'h5; //< 
    18'h16622: Data = 4'h5; //< 
    18'h16623: Data = 4'h6; //[ 
    18'h16624: Data = 4'h3; //- 
    18'h16625: Data = 4'h4; //> 
    18'h16626: Data = 4'h4; //> 
    18'h16627: Data = 4'h4; //> 
    18'h16628: Data = 4'h3; //- 
    18'h16629: Data = 4'h5; //< 
    18'h16630: Data = 4'h5; //< 
    18'h16631: Data = 4'h5; //< 
    18'h16632: Data = 4'h5; //< 
    18'h16633: Data = 4'h5; //< 
    18'h16634: Data = 4'h5; //< 
    18'h16635: Data = 4'h5; //< 
    18'h16636: Data = 4'h5; //< 
    18'h16637: Data = 4'h5; //< 
    18'h16638: Data = 4'h5; //< 
    18'h16639: Data = 4'h5; //< 
    18'h16640: Data = 4'h5; //< 
    18'h16641: Data = 4'h5; //< 
    18'h16642: Data = 4'h2; //+ 
    18'h16643: Data = 4'h4; //> 
    18'h16644: Data = 4'h4; //> 
    18'h16645: Data = 4'h4; //> 
    18'h16646: Data = 4'h4; //> 
    18'h16647: Data = 4'h4; //> 
    18'h16648: Data = 4'h4; //> 
    18'h16649: Data = 4'h4; //> 
    18'h16650: Data = 4'h4; //> 
    18'h16651: Data = 4'h4; //> 
    18'h16652: Data = 4'h4; //> 
    18'h16653: Data = 4'h7; //] 
    18'h16654: Data = 4'h4; //> 
    18'h16655: Data = 4'h7; //] 
    18'h16656: Data = 4'h5; //< 
    18'h16657: Data = 4'h6; //[ 
    18'h16658: Data = 4'h3; //- 
    18'h16659: Data = 4'h4; //> 
    18'h16660: Data = 4'h4; //> 
    18'h16661: Data = 4'h4; //> 
    18'h16662: Data = 4'h2; //+ 
    18'h16663: Data = 4'h5; //< 
    18'h16664: Data = 4'h5; //< 
    18'h16665: Data = 4'h5; //< 
    18'h16666: Data = 4'h7; //] 
    18'h16667: Data = 4'h5; //< 
    18'h16668: Data = 4'h5; //< 
    18'h16669: Data = 4'h5; //< 
    18'h16670: Data = 4'h5; //< 
    18'h16671: Data = 4'h5; //< 
    18'h16672: Data = 4'h5; //< 
    18'h16673: Data = 4'h5; //< 
    18'h16674: Data = 4'h5; //< 
    18'h16675: Data = 4'h5; //< 
    18'h16676: Data = 4'h5; //< 
    18'h16677: Data = 4'h5; //< 
    18'h16678: Data = 4'h7; //] 
    18'h16679: Data = 4'h4; //> 
    18'h16680: Data = 4'h4; //> 
    18'h16681: Data = 4'h4; //> 
    18'h16682: Data = 4'h4; //> 
    18'h16683: Data = 4'h4; //> 
    18'h16684: Data = 4'ha; //0 
    18'h16685: Data = 4'h4; //> 
    18'h16686: Data = 4'h4; //> 
    18'h16687: Data = 4'h6; //[ 
    18'h16688: Data = 4'h3; //- 
    18'h16689: Data = 4'h5; //< 
    18'h16690: Data = 4'h5; //< 
    18'h16691: Data = 4'h5; //< 
    18'h16692: Data = 4'h5; //< 
    18'h16693: Data = 4'h5; //< 
    18'h16694: Data = 4'h5; //< 
    18'h16695: Data = 4'h5; //< 
    18'h16696: Data = 4'h2; //+ 
    18'h16697: Data = 4'h4; //> 
    18'h16698: Data = 4'h4; //> 
    18'h16699: Data = 4'h4; //> 
    18'h16700: Data = 4'h4; //> 
    18'h16701: Data = 4'h4; //> 
    18'h16702: Data = 4'h4; //> 
    18'h16703: Data = 4'h4; //> 
    18'h16704: Data = 4'h7; //] 
    18'h16705: Data = 4'h5; //< 
    18'h16706: Data = 4'h5; //< 
    18'h16707: Data = 4'h5; //< 
    18'h16708: Data = 4'h5; //< 
    18'h16709: Data = 4'h5; //< 
    18'h16710: Data = 4'h5; //< 
    18'h16711: Data = 4'h5; //< 
    18'h16712: Data = 4'h6; //[ 
    18'h16713: Data = 4'h3; //- 
    18'h16714: Data = 4'h4; //> 
    18'h16715: Data = 4'h4; //> 
    18'h16716: Data = 4'h4; //> 
    18'h16717: Data = 4'h4; //> 
    18'h16718: Data = 4'h4; //> 
    18'h16719: Data = 4'h4; //> 
    18'h16720: Data = 4'h4; //> 
    18'h16721: Data = 4'h2; //+ 
    18'h16722: Data = 4'h5; //< 
    18'h16723: Data = 4'h5; //< 
    18'h16724: Data = 4'h2; //+ 
    18'h16725: Data = 4'h5; //< 
    18'h16726: Data = 4'h5; //< 
    18'h16727: Data = 4'h5; //< 
    18'h16728: Data = 4'h5; //< 
    18'h16729: Data = 4'h5; //< 
    18'h16730: Data = 4'h7; //] 
    18'h16731: Data = 4'h7; //] 
    18'h16732: Data = 4'h4; //> 
    18'h16733: Data = 4'h4; //> 
    18'h16734: Data = 4'h4; //> 
    18'h16735: Data = 4'h4; //> 
    18'h16736: Data = 4'h6; //[ 
    18'h16737: Data = 4'h3; //- 
    18'h16738: Data = 4'h5; //< 
    18'h16739: Data = 4'h5; //< 
    18'h16740: Data = 4'h5; //< 
    18'h16741: Data = 4'h5; //< 
    18'h16742: Data = 4'h2; //+ 
    18'h16743: Data = 4'h4; //> 
    18'h16744: Data = 4'h4; //> 
    18'h16745: Data = 4'h4; //> 
    18'h16746: Data = 4'h4; //> 
    18'h16747: Data = 4'h7; //] 
    18'h16748: Data = 4'h5; //< 
    18'h16749: Data = 4'h5; //< 
    18'h16750: Data = 4'h5; //< 
    18'h16751: Data = 4'h5; //< 
    18'h16752: Data = 4'h6; //[ 
    18'h16753: Data = 4'h3; //- 
    18'h16754: Data = 4'h4; //> 
    18'h16755: Data = 4'h4; //> 
    18'h16756: Data = 4'h4; //> 
    18'h16757: Data = 4'h4; //> 
    18'h16758: Data = 4'h2; //+ 
    18'h16759: Data = 4'h4; //> 
    18'h16760: Data = 4'h4; //> 
    18'h16761: Data = 4'h4; //> 
    18'h16762: Data = 4'h4; //> 
    18'h16763: Data = 4'h4; //> 
    18'h16764: Data = 4'h6; //[ 
    18'h16765: Data = 4'h4; //> 
    18'h16766: Data = 4'h2; //+ 
    18'h16767: Data = 4'h4; //> 
    18'h16768: Data = 4'h4; //> 
    18'h16769: Data = 4'h6; //[ 
    18'h16770: Data = 4'h3; //- 
    18'h16771: Data = 4'h5; //< 
    18'h16772: Data = 4'h5; //< 
    18'h16773: Data = 4'h3; //- 
    18'h16774: Data = 4'h4; //> 
    18'h16775: Data = 4'h4; //> 
    18'h16776: Data = 4'h7; //] 
    18'h16777: Data = 4'h5; //< 
    18'h16778: Data = 4'h5; //< 
    18'h16779: Data = 4'h6; //[ 
    18'h16780: Data = 4'h3; //- 
    18'h16781: Data = 4'h4; //> 
    18'h16782: Data = 4'h4; //> 
    18'h16783: Data = 4'h2; //+ 
    18'h16784: Data = 4'h5; //< 
    18'h16785: Data = 4'h5; //< 
    18'h16786: Data = 4'h7; //] 
    18'h16787: Data = 4'h4; //> 
    18'h16788: Data = 4'h4; //> 
    18'h16789: Data = 4'h4; //> 
    18'h16790: Data = 4'h4; //> 
    18'h16791: Data = 4'h4; //> 
    18'h16792: Data = 4'h4; //> 
    18'h16793: Data = 4'h4; //> 
    18'h16794: Data = 4'h4; //> 
    18'h16795: Data = 4'h7; //] 
    18'h16796: Data = 4'h5; //< 
    18'h16797: Data = 4'h5; //< 
    18'h16798: Data = 4'h5; //< 
    18'h16799: Data = 4'h5; //< 
    18'h16800: Data = 4'h5; //< 
    18'h16801: Data = 4'h5; //< 
    18'h16802: Data = 4'h5; //< 
    18'h16803: Data = 4'h5; //< 
    18'h16804: Data = 4'h2; //+ 
    18'h16805: Data = 4'h5; //< 
    18'h16806: Data = 4'h6; //[ 
    18'h16807: Data = 4'h4; //> 
    18'h16808: Data = 4'h6; //[ 
    18'h16809: Data = 4'h3; //- 
    18'h16810: Data = 4'h4; //> 
    18'h16811: Data = 4'h4; //> 
    18'h16812: Data = 4'h4; //> 
    18'h16813: Data = 4'h4; //> 
    18'h16814: Data = 4'h2; //+ 
    18'h16815: Data = 4'h5; //< 
    18'h16816: Data = 4'h5; //< 
    18'h16817: Data = 4'h5; //< 
    18'h16818: Data = 4'h6; //[ 
    18'h16819: Data = 4'h3; //- 
    18'h16820: Data = 4'h4; //> 
    18'h16821: Data = 4'h4; //> 
    18'h16822: Data = 4'h4; //> 
    18'h16823: Data = 4'h3; //- 
    18'h16824: Data = 4'h5; //< 
    18'h16825: Data = 4'h5; //< 
    18'h16826: Data = 4'h5; //< 
    18'h16827: Data = 4'h5; //< 
    18'h16828: Data = 4'h5; //< 
    18'h16829: Data = 4'h5; //< 
    18'h16830: Data = 4'h5; //< 
    18'h16831: Data = 4'h5; //< 
    18'h16832: Data = 4'h5; //< 
    18'h16833: Data = 4'h5; //< 
    18'h16834: Data = 4'h5; //< 
    18'h16835: Data = 4'h5; //< 
    18'h16836: Data = 4'h5; //< 
    18'h16837: Data = 4'h2; //+ 
    18'h16838: Data = 4'h4; //> 
    18'h16839: Data = 4'h4; //> 
    18'h16840: Data = 4'h4; //> 
    18'h16841: Data = 4'h4; //> 
    18'h16842: Data = 4'h4; //> 
    18'h16843: Data = 4'h4; //> 
    18'h16844: Data = 4'h4; //> 
    18'h16845: Data = 4'h4; //> 
    18'h16846: Data = 4'h4; //> 
    18'h16847: Data = 4'h4; //> 
    18'h16848: Data = 4'h4; //> 
    18'h16849: Data = 4'h6; //[ 
    18'h16850: Data = 4'h3; //- 
    18'h16851: Data = 4'h4; //> 
    18'h16852: Data = 4'h4; //> 
    18'h16853: Data = 4'h2; //+ 
    18'h16854: Data = 4'h5; //< 
    18'h16855: Data = 4'h5; //< 
    18'h16856: Data = 4'h7; //] 
    18'h16857: Data = 4'h5; //< 
    18'h16858: Data = 4'h7; //] 
    18'h16859: Data = 4'h4; //> 
    18'h16860: Data = 4'h6; //[ 
    18'h16861: Data = 4'h3; //- 
    18'h16862: Data = 4'h4; //> 
    18'h16863: Data = 4'h4; //> 
    18'h16864: Data = 4'h3; //- 
    18'h16865: Data = 4'h5; //< 
    18'h16866: Data = 4'h5; //< 
    18'h16867: Data = 4'h5; //< 
    18'h16868: Data = 4'h5; //< 
    18'h16869: Data = 4'h5; //< 
    18'h16870: Data = 4'h5; //< 
    18'h16871: Data = 4'h5; //< 
    18'h16872: Data = 4'h5; //< 
    18'h16873: Data = 4'h5; //< 
    18'h16874: Data = 4'h5; //< 
    18'h16875: Data = 4'h5; //< 
    18'h16876: Data = 4'h5; //< 
    18'h16877: Data = 4'h5; //< 
    18'h16878: Data = 4'h2; //+ 
    18'h16879: Data = 4'h4; //> 
    18'h16880: Data = 4'h4; //> 
    18'h16881: Data = 4'h4; //> 
    18'h16882: Data = 4'h4; //> 
    18'h16883: Data = 4'h4; //> 
    18'h16884: Data = 4'h4; //> 
    18'h16885: Data = 4'h4; //> 
    18'h16886: Data = 4'h4; //> 
    18'h16887: Data = 4'h4; //> 
    18'h16888: Data = 4'h4; //> 
    18'h16889: Data = 4'h4; //> 
    18'h16890: Data = 4'h7; //] 
    18'h16891: Data = 4'h5; //< 
    18'h16892: Data = 4'h5; //< 
    18'h16893: Data = 4'h7; //] 
    18'h16894: Data = 4'h4; //> 
    18'h16895: Data = 4'h6; //[ 
    18'h16896: Data = 4'h3; //- 
    18'h16897: Data = 4'h4; //> 
    18'h16898: Data = 4'h4; //> 
    18'h16899: Data = 4'h4; //> 
    18'h16900: Data = 4'h2; //+ 
    18'h16901: Data = 4'h5; //< 
    18'h16902: Data = 4'h5; //< 
    18'h16903: Data = 4'h6; //[ 
    18'h16904: Data = 4'h3; //- 
    18'h16905: Data = 4'h4; //> 
    18'h16906: Data = 4'h4; //> 
    18'h16907: Data = 4'h3; //- 
    18'h16908: Data = 4'h5; //< 
    18'h16909: Data = 4'h5; //< 
    18'h16910: Data = 4'h5; //< 
    18'h16911: Data = 4'h5; //< 
    18'h16912: Data = 4'h5; //< 
    18'h16913: Data = 4'h5; //< 
    18'h16914: Data = 4'h5; //< 
    18'h16915: Data = 4'h5; //< 
    18'h16916: Data = 4'h5; //< 
    18'h16917: Data = 4'h5; //< 
    18'h16918: Data = 4'h5; //< 
    18'h16919: Data = 4'h5; //< 
    18'h16920: Data = 4'h5; //< 
    18'h16921: Data = 4'h2; //+ 
    18'h16922: Data = 4'h4; //> 
    18'h16923: Data = 4'h4; //> 
    18'h16924: Data = 4'h4; //> 
    18'h16925: Data = 4'h4; //> 
    18'h16926: Data = 4'h4; //> 
    18'h16927: Data = 4'h4; //> 
    18'h16928: Data = 4'h4; //> 
    18'h16929: Data = 4'h4; //> 
    18'h16930: Data = 4'h4; //> 
    18'h16931: Data = 4'h4; //> 
    18'h16932: Data = 4'h4; //> 
    18'h16933: Data = 4'h7; //] 
    18'h16934: Data = 4'h5; //< 
    18'h16935: Data = 4'h7; //] 
    18'h16936: Data = 4'h4; //> 
    18'h16937: Data = 4'h6; //[ 
    18'h16938: Data = 4'h3; //- 
    18'h16939: Data = 4'h4; //> 
    18'h16940: Data = 4'h4; //> 
    18'h16941: Data = 4'h2; //+ 
    18'h16942: Data = 4'h5; //< 
    18'h16943: Data = 4'h5; //< 
    18'h16944: Data = 4'h7; //] 
    18'h16945: Data = 4'h5; //< 
    18'h16946: Data = 4'h5; //< 
    18'h16947: Data = 4'h5; //< 
    18'h16948: Data = 4'h5; //< 
    18'h16949: Data = 4'h5; //< 
    18'h16950: Data = 4'h5; //< 
    18'h16951: Data = 4'h5; //< 
    18'h16952: Data = 4'h5; //< 
    18'h16953: Data = 4'h5; //< 
    18'h16954: Data = 4'h5; //< 
    18'h16955: Data = 4'h5; //< 
    18'h16956: Data = 4'h5; //< 
    18'h16957: Data = 4'h7; //] 
    18'h16958: Data = 4'h7; //] 
    18'h16959: Data = 4'h4; //> 
    18'h16960: Data = 4'h4; //> 
    18'h16961: Data = 4'h4; //> 
    18'h16962: Data = 4'h4; //> 
    18'h16963: Data = 4'ha; //0 
    18'h16964: Data = 4'h5; //< 
    18'h16965: Data = 4'h5; //< 
    18'h16966: Data = 4'h5; //< 
    18'h16967: Data = 4'h5; //< 
    18'h16968: Data = 4'h7; //] 
    18'h16969: Data = 4'h4; //> 
    18'h16970: Data = 4'h4; //> 
    18'h16971: Data = 4'h4; //> 
    18'h16972: Data = 4'h4; //> 
    18'h16973: Data = 4'h6; //[ 
    18'h16974: Data = 4'h3; //- 
    18'h16975: Data = 4'h5; //< 
    18'h16976: Data = 4'h5; //< 
    18'h16977: Data = 4'h5; //< 
    18'h16978: Data = 4'h5; //< 
    18'h16979: Data = 4'h2; //+ 
    18'h16980: Data = 4'h4; //> 
    18'h16981: Data = 4'h4; //> 
    18'h16982: Data = 4'h4; //> 
    18'h16983: Data = 4'h4; //> 
    18'h16984: Data = 4'h7; //] 
    18'h16985: Data = 4'h5; //< 
    18'h16986: Data = 4'h5; //< 
    18'h16987: Data = 4'h5; //< 
    18'h16988: Data = 4'h5; //< 
    18'h16989: Data = 4'h6; //[ 
    18'h16990: Data = 4'h3; //- 
    18'h16991: Data = 4'h4; //> 
    18'h16992: Data = 4'h4; //> 
    18'h16993: Data = 4'h4; //> 
    18'h16994: Data = 4'h4; //> 
    18'h16995: Data = 4'h2; //+ 
    18'h16996: Data = 4'h4; //> 
    18'h16997: Data = 4'ha; //0 
    18'h16998: Data = 4'h4; //> 
    18'h16999: Data = 4'h4; //> 
    18'h17000: Data = 4'h6; //[ 
    18'h17001: Data = 4'h3; //- 
    18'h17002: Data = 4'h5; //< 
    18'h17003: Data = 4'h5; //< 
    18'h17004: Data = 4'h5; //< 
    18'h17005: Data = 4'h5; //< 
    18'h17006: Data = 4'h5; //< 
    18'h17007: Data = 4'h5; //< 
    18'h17008: Data = 4'h5; //< 
    18'h17009: Data = 4'h2; //+ 
    18'h17010: Data = 4'h4; //> 
    18'h17011: Data = 4'h4; //> 
    18'h17012: Data = 4'h4; //> 
    18'h17013: Data = 4'h4; //> 
    18'h17014: Data = 4'h4; //> 
    18'h17015: Data = 4'h4; //> 
    18'h17016: Data = 4'h4; //> 
    18'h17017: Data = 4'h7; //] 
    18'h17018: Data = 4'h5; //< 
    18'h17019: Data = 4'h5; //< 
    18'h17020: Data = 4'h5; //< 
    18'h17021: Data = 4'h5; //< 
    18'h17022: Data = 4'h5; //< 
    18'h17023: Data = 4'h5; //< 
    18'h17024: Data = 4'h5; //< 
    18'h17025: Data = 4'h6; //[ 
    18'h17026: Data = 4'h3; //- 
    18'h17027: Data = 4'h4; //> 
    18'h17028: Data = 4'h4; //> 
    18'h17029: Data = 4'h4; //> 
    18'h17030: Data = 4'h4; //> 
    18'h17031: Data = 4'h4; //> 
    18'h17032: Data = 4'h4; //> 
    18'h17033: Data = 4'h4; //> 
    18'h17034: Data = 4'h2; //+ 
    18'h17035: Data = 4'h5; //< 
    18'h17036: Data = 4'h5; //< 
    18'h17037: Data = 4'h2; //+ 
    18'h17038: Data = 4'h5; //< 
    18'h17039: Data = 4'h5; //< 
    18'h17040: Data = 4'h5; //< 
    18'h17041: Data = 4'h5; //< 
    18'h17042: Data = 4'h5; //< 
    18'h17043: Data = 4'h7; //] 
    18'h17044: Data = 4'h4; //> 
    18'h17045: Data = 4'h4; //> 
    18'h17046: Data = 4'h4; //> 
    18'h17047: Data = 4'h4; //> 
    18'h17048: Data = 4'h4; //> 
    18'h17049: Data = 4'h4; //> 
    18'h17050: Data = 4'h4; //> 
    18'h17051: Data = 4'h4; //> 
    18'h17052: Data = 4'h4; //> 
    18'h17053: Data = 4'h6; //[ 
    18'h17054: Data = 4'h4; //> 
    18'h17055: Data = 4'h4; //> 
    18'h17056: Data = 4'h4; //> 
    18'h17057: Data = 4'h4; //> 
    18'h17058: Data = 4'h4; //> 
    18'h17059: Data = 4'h4; //> 
    18'h17060: Data = 4'h4; //> 
    18'h17061: Data = 4'h4; //> 
    18'h17062: Data = 4'h4; //> 
    18'h17063: Data = 4'h7; //] 
    18'h17064: Data = 4'h5; //< 
    18'h17065: Data = 4'h5; //< 
    18'h17066: Data = 4'h5; //< 
    18'h17067: Data = 4'h5; //< 
    18'h17068: Data = 4'h5; //< 
    18'h17069: Data = 4'h5; //< 
    18'h17070: Data = 4'h5; //< 
    18'h17071: Data = 4'h5; //< 
    18'h17072: Data = 4'h5; //< 
    18'h17073: Data = 4'h6; //[ 
    18'h17074: Data = 4'h4; //> 
    18'h17075: Data = 4'h6; //[ 
    18'h17076: Data = 4'h3; //- 
    18'h17077: Data = 4'h4; //> 
    18'h17078: Data = 4'h4; //> 
    18'h17079: Data = 4'h4; //> 
    18'h17080: Data = 4'h4; //> 
    18'h17081: Data = 4'h2; //+ 
    18'h17082: Data = 4'h5; //< 
    18'h17083: Data = 4'h5; //< 
    18'h17084: Data = 4'h5; //< 
    18'h17085: Data = 4'h6; //[ 
    18'h17086: Data = 4'h3; //- 
    18'h17087: Data = 4'h4; //> 
    18'h17088: Data = 4'h4; //> 
    18'h17089: Data = 4'h4; //> 
    18'h17090: Data = 4'h3; //- 
    18'h17091: Data = 4'h5; //< 
    18'h17092: Data = 4'h5; //< 
    18'h17093: Data = 4'h5; //< 
    18'h17094: Data = 4'h5; //< 
    18'h17095: Data = 4'h5; //< 
    18'h17096: Data = 4'h5; //< 
    18'h17097: Data = 4'h5; //< 
    18'h17098: Data = 4'h5; //< 
    18'h17099: Data = 4'h5; //< 
    18'h17100: Data = 4'h5; //< 
    18'h17101: Data = 4'h5; //< 
    18'h17102: Data = 4'h5; //< 
    18'h17103: Data = 4'h5; //< 
    18'h17104: Data = 4'h2; //+ 
    18'h17105: Data = 4'h4; //> 
    18'h17106: Data = 4'h4; //> 
    18'h17107: Data = 4'h4; //> 
    18'h17108: Data = 4'h4; //> 
    18'h17109: Data = 4'h4; //> 
    18'h17110: Data = 4'h4; //> 
    18'h17111: Data = 4'h4; //> 
    18'h17112: Data = 4'h4; //> 
    18'h17113: Data = 4'h4; //> 
    18'h17114: Data = 4'h4; //> 
    18'h17115: Data = 4'h4; //> 
    18'h17116: Data = 4'h6; //[ 
    18'h17117: Data = 4'h3; //- 
    18'h17118: Data = 4'h4; //> 
    18'h17119: Data = 4'h4; //> 
    18'h17120: Data = 4'h2; //+ 
    18'h17121: Data = 4'h5; //< 
    18'h17122: Data = 4'h5; //< 
    18'h17123: Data = 4'h7; //] 
    18'h17124: Data = 4'h5; //< 
    18'h17125: Data = 4'h7; //] 
    18'h17126: Data = 4'h4; //> 
    18'h17127: Data = 4'h6; //[ 
    18'h17128: Data = 4'h3; //- 
    18'h17129: Data = 4'h4; //> 
    18'h17130: Data = 4'h4; //> 
    18'h17131: Data = 4'h3; //- 
    18'h17132: Data = 4'h5; //< 
    18'h17133: Data = 4'h5; //< 
    18'h17134: Data = 4'h5; //< 
    18'h17135: Data = 4'h5; //< 
    18'h17136: Data = 4'h5; //< 
    18'h17137: Data = 4'h5; //< 
    18'h17138: Data = 4'h5; //< 
    18'h17139: Data = 4'h5; //< 
    18'h17140: Data = 4'h5; //< 
    18'h17141: Data = 4'h5; //< 
    18'h17142: Data = 4'h5; //< 
    18'h17143: Data = 4'h5; //< 
    18'h17144: Data = 4'h5; //< 
    18'h17145: Data = 4'h2; //+ 
    18'h17146: Data = 4'h4; //> 
    18'h17147: Data = 4'h4; //> 
    18'h17148: Data = 4'h4; //> 
    18'h17149: Data = 4'h4; //> 
    18'h17150: Data = 4'h4; //> 
    18'h17151: Data = 4'h4; //> 
    18'h17152: Data = 4'h4; //> 
    18'h17153: Data = 4'h4; //> 
    18'h17154: Data = 4'h4; //> 
    18'h17155: Data = 4'h4; //> 
    18'h17156: Data = 4'h4; //> 
    18'h17157: Data = 4'h7; //] 
    18'h17158: Data = 4'h5; //< 
    18'h17159: Data = 4'h5; //< 
    18'h17160: Data = 4'h7; //] 
    18'h17161: Data = 4'h4; //> 
    18'h17162: Data = 4'h6; //[ 
    18'h17163: Data = 4'h3; //- 
    18'h17164: Data = 4'h4; //> 
    18'h17165: Data = 4'h4; //> 
    18'h17166: Data = 4'h4; //> 
    18'h17167: Data = 4'h2; //+ 
    18'h17168: Data = 4'h5; //< 
    18'h17169: Data = 4'h5; //< 
    18'h17170: Data = 4'h6; //[ 
    18'h17171: Data = 4'h3; //- 
    18'h17172: Data = 4'h4; //> 
    18'h17173: Data = 4'h4; //> 
    18'h17174: Data = 4'h3; //- 
    18'h17175: Data = 4'h5; //< 
    18'h17176: Data = 4'h5; //< 
    18'h17177: Data = 4'h5; //< 
    18'h17178: Data = 4'h5; //< 
    18'h17179: Data = 4'h5; //< 
    18'h17180: Data = 4'h5; //< 
    18'h17181: Data = 4'h5; //< 
    18'h17182: Data = 4'h5; //< 
    18'h17183: Data = 4'h5; //< 
    18'h17184: Data = 4'h5; //< 
    18'h17185: Data = 4'h5; //< 
    18'h17186: Data = 4'h5; //< 
    18'h17187: Data = 4'h5; //< 
    18'h17188: Data = 4'h2; //+ 
    18'h17189: Data = 4'h4; //> 
    18'h17190: Data = 4'h4; //> 
    18'h17191: Data = 4'h4; //> 
    18'h17192: Data = 4'h4; //> 
    18'h17193: Data = 4'h4; //> 
    18'h17194: Data = 4'h4; //> 
    18'h17195: Data = 4'h4; //> 
    18'h17196: Data = 4'h4; //> 
    18'h17197: Data = 4'h4; //> 
    18'h17198: Data = 4'h4; //> 
    18'h17199: Data = 4'h4; //> 
    18'h17200: Data = 4'h7; //] 
    18'h17201: Data = 4'h5; //< 
    18'h17202: Data = 4'h7; //] 
    18'h17203: Data = 4'h4; //> 
    18'h17204: Data = 4'h6; //[ 
    18'h17205: Data = 4'h3; //- 
    18'h17206: Data = 4'h4; //> 
    18'h17207: Data = 4'h4; //> 
    18'h17208: Data = 4'h2; //+ 
    18'h17209: Data = 4'h5; //< 
    18'h17210: Data = 4'h5; //< 
    18'h17211: Data = 4'h7; //] 
    18'h17212: Data = 4'h5; //< 
    18'h17213: Data = 4'h5; //< 
    18'h17214: Data = 4'h5; //< 
    18'h17215: Data = 4'h5; //< 
    18'h17216: Data = 4'h5; //< 
    18'h17217: Data = 4'h5; //< 
    18'h17218: Data = 4'h5; //< 
    18'h17219: Data = 4'h5; //< 
    18'h17220: Data = 4'h5; //< 
    18'h17221: Data = 4'h5; //< 
    18'h17222: Data = 4'h5; //< 
    18'h17223: Data = 4'h5; //< 
    18'h17224: Data = 4'h7; //] 
    18'h17225: Data = 4'h7; //] 
    18'h17226: Data = 4'h4; //> 
    18'h17227: Data = 4'h4; //> 
    18'h17228: Data = 4'h4; //> 
    18'h17229: Data = 4'h4; //> 
    18'h17230: Data = 4'h4; //> 
    18'h17231: Data = 4'h4; //> 
    18'h17232: Data = 4'h4; //> 
    18'h17233: Data = 4'h4; //> 
    18'h17234: Data = 4'h4; //> 
    18'h17235: Data = 4'h6; //[ 
    18'h17236: Data = 4'h4; //> 
    18'h17237: Data = 4'h4; //> 
    18'h17238: Data = 4'ha; //0 
    18'h17239: Data = 4'h4; //> 
    18'h17240: Data = 4'ha; //0 
    18'h17241: Data = 4'h4; //> 
    18'h17242: Data = 4'h4; //> 
    18'h17243: Data = 4'h4; //> 
    18'h17244: Data = 4'h4; //> 
    18'h17245: Data = 4'h4; //> 
    18'h17246: Data = 4'h4; //> 
    18'h17247: Data = 4'h7; //] 
    18'h17248: Data = 4'h5; //< 
    18'h17249: Data = 4'h5; //< 
    18'h17250: Data = 4'h5; //< 
    18'h17251: Data = 4'h5; //< 
    18'h17252: Data = 4'h5; //< 
    18'h17253: Data = 4'h5; //< 
    18'h17254: Data = 4'h5; //< 
    18'h17255: Data = 4'h5; //< 
    18'h17256: Data = 4'h5; //< 
    18'h17257: Data = 4'h6; //[ 
    18'h17258: Data = 4'h5; //< 
    18'h17259: Data = 4'h5; //< 
    18'h17260: Data = 4'h5; //< 
    18'h17261: Data = 4'h5; //< 
    18'h17262: Data = 4'h5; //< 
    18'h17263: Data = 4'h5; //< 
    18'h17264: Data = 4'h5; //< 
    18'h17265: Data = 4'h5; //< 
    18'h17266: Data = 4'h5; //< 
    18'h17267: Data = 4'h7; //] 
    18'h17268: Data = 4'h4; //> 
    18'h17269: Data = 4'h4; //> 
    18'h17270: Data = 4'h4; //> 
    18'h17271: Data = 4'ha; //0 
    18'h17272: Data = 4'h4; //> 
    18'h17273: Data = 4'ha; //0 
    18'h17274: Data = 4'h4; //> 
    18'h17275: Data = 4'h4; //> 
    18'h17276: Data = 4'h4; //> 
    18'h17277: Data = 4'h4; //> 
    18'h17278: Data = 4'h4; //> 
    18'h17279: Data = 4'h6; //[ 
    18'h17280: Data = 4'h4; //> 
    18'h17281: Data = 4'h4; //> 
    18'h17282: Data = 4'h4; //> 
    18'h17283: Data = 4'h4; //> 
    18'h17284: Data = 4'h4; //> 
    18'h17285: Data = 4'h6; //[ 
    18'h17286: Data = 4'h3; //- 
    18'h17287: Data = 4'h5; //< 
    18'h17288: Data = 4'h5; //< 
    18'h17289: Data = 4'h5; //< 
    18'h17290: Data = 4'h5; //< 
    18'h17291: Data = 4'h2; //+ 
    18'h17292: Data = 4'h4; //> 
    18'h17293: Data = 4'h4; //> 
    18'h17294: Data = 4'h4; //> 
    18'h17295: Data = 4'h4; //> 
    18'h17296: Data = 4'h7; //] 
    18'h17297: Data = 4'h5; //< 
    18'h17298: Data = 4'h5; //< 
    18'h17299: Data = 4'h5; //< 
    18'h17300: Data = 4'h5; //< 
    18'h17301: Data = 4'h6; //[ 
    18'h17302: Data = 4'h3; //- 
    18'h17303: Data = 4'h4; //> 
    18'h17304: Data = 4'h4; //> 
    18'h17305: Data = 4'h4; //> 
    18'h17306: Data = 4'h4; //> 
    18'h17307: Data = 4'h2; //+ 
    18'h17308: Data = 4'h5; //< 
    18'h17309: Data = 4'h5; //< 
    18'h17310: Data = 4'h5; //< 
    18'h17311: Data = 4'h2; //+ 
    18'h17312: Data = 4'h5; //< 
    18'h17313: Data = 4'h7; //] 
    18'h17314: Data = 4'h4; //> 
    18'h17315: Data = 4'h4; //> 
    18'h17316: Data = 4'h4; //> 
    18'h17317: Data = 4'h4; //> 
    18'h17318: Data = 4'h4; //> 
    18'h17319: Data = 4'h4; //> 
    18'h17320: Data = 4'h4; //> 
    18'h17321: Data = 4'h4; //> 
    18'h17322: Data = 4'h7; //] 
    18'h17323: Data = 4'h5; //< 
    18'h17324: Data = 4'h5; //< 
    18'h17325: Data = 4'h5; //< 
    18'h17326: Data = 4'h5; //< 
    18'h17327: Data = 4'h5; //< 
    18'h17328: Data = 4'h5; //< 
    18'h17329: Data = 4'h5; //< 
    18'h17330: Data = 4'h5; //< 
    18'h17331: Data = 4'h5; //< 
    18'h17332: Data = 4'h6; //[ 
    18'h17333: Data = 4'h5; //< 
    18'h17334: Data = 4'h5; //< 
    18'h17335: Data = 4'h5; //< 
    18'h17336: Data = 4'h5; //< 
    18'h17337: Data = 4'h5; //< 
    18'h17338: Data = 4'h5; //< 
    18'h17339: Data = 4'h5; //< 
    18'h17340: Data = 4'h5; //< 
    18'h17341: Data = 4'h5; //< 
    18'h17342: Data = 4'h7; //] 
    18'h17343: Data = 4'h4; //> 
    18'h17344: Data = 4'h4; //> 
    18'h17345: Data = 4'h4; //> 
    18'h17346: Data = 4'h4; //> 
    18'h17347: Data = 4'h4; //> 
    18'h17348: Data = 4'h4; //> 
    18'h17349: Data = 4'h4; //> 
    18'h17350: Data = 4'h4; //> 
    18'h17351: Data = 4'h4; //> 
    18'h17352: Data = 4'h6; //[ 
    18'h17353: Data = 4'h4; //> 
    18'h17354: Data = 4'h4; //> 
    18'h17355: Data = 4'h4; //> 
    18'h17356: Data = 4'h4; //> 
    18'h17357: Data = 4'h4; //> 
    18'h17358: Data = 4'h4; //> 
    18'h17359: Data = 4'h6; //[ 
    18'h17360: Data = 4'h3; //- 
    18'h17361: Data = 4'h5; //< 
    18'h17362: Data = 4'h5; //< 
    18'h17363: Data = 4'h5; //< 
    18'h17364: Data = 4'h5; //< 
    18'h17365: Data = 4'h5; //< 
    18'h17366: Data = 4'h2; //+ 
    18'h17367: Data = 4'h4; //> 
    18'h17368: Data = 4'h4; //> 
    18'h17369: Data = 4'h4; //> 
    18'h17370: Data = 4'h4; //> 
    18'h17371: Data = 4'h4; //> 
    18'h17372: Data = 4'h7; //] 
    18'h17373: Data = 4'h5; //< 
    18'h17374: Data = 4'h5; //< 
    18'h17375: Data = 4'h5; //< 
    18'h17376: Data = 4'h5; //< 
    18'h17377: Data = 4'h5; //< 
    18'h17378: Data = 4'h6; //[ 
    18'h17379: Data = 4'h3; //- 
    18'h17380: Data = 4'h4; //> 
    18'h17381: Data = 4'h4; //> 
    18'h17382: Data = 4'h4; //> 
    18'h17383: Data = 4'h4; //> 
    18'h17384: Data = 4'h4; //> 
    18'h17385: Data = 4'h2; //+ 
    18'h17386: Data = 4'h5; //< 
    18'h17387: Data = 4'h5; //< 
    18'h17388: Data = 4'h5; //< 
    18'h17389: Data = 4'h2; //+ 
    18'h17390: Data = 4'h5; //< 
    18'h17391: Data = 4'h5; //< 
    18'h17392: Data = 4'h7; //] 
    18'h17393: Data = 4'h4; //> 
    18'h17394: Data = 4'h4; //> 
    18'h17395: Data = 4'h4; //> 
    18'h17396: Data = 4'h4; //> 
    18'h17397: Data = 4'h4; //> 
    18'h17398: Data = 4'h4; //> 
    18'h17399: Data = 4'h4; //> 
    18'h17400: Data = 4'h4; //> 
    18'h17401: Data = 4'h7; //] 
    18'h17402: Data = 4'h5; //< 
    18'h17403: Data = 4'h5; //< 
    18'h17404: Data = 4'h5; //< 
    18'h17405: Data = 4'h5; //< 
    18'h17406: Data = 4'h5; //< 
    18'h17407: Data = 4'h5; //< 
    18'h17408: Data = 4'h5; //< 
    18'h17409: Data = 4'h5; //< 
    18'h17410: Data = 4'h5; //< 
    18'h17411: Data = 4'h6; //[ 
    18'h17412: Data = 4'h5; //< 
    18'h17413: Data = 4'h5; //< 
    18'h17414: Data = 4'h5; //< 
    18'h17415: Data = 4'h5; //< 
    18'h17416: Data = 4'h5; //< 
    18'h17417: Data = 4'h5; //< 
    18'h17418: Data = 4'h5; //< 
    18'h17419: Data = 4'h5; //< 
    18'h17420: Data = 4'h5; //< 
    18'h17421: Data = 4'h7; //] 
    18'h17422: Data = 4'h4; //> 
    18'h17423: Data = 4'h4; //> 
    18'h17424: Data = 4'h4; //> 
    18'h17425: Data = 4'h4; //> 
    18'h17426: Data = 4'h4; //> 
    18'h17427: Data = 4'h4; //> 
    18'h17428: Data = 4'h4; //> 
    18'h17429: Data = 4'h4; //> 
    18'h17430: Data = 4'h4; //> 
    18'h17431: Data = 4'h2; //+ 
    18'h17432: Data = 4'h2; //+ 
    18'h17433: Data = 4'h2; //+ 
    18'h17434: Data = 4'h2; //+ 
    18'h17435: Data = 4'h2; //+ 
    18'h17436: Data = 4'h2; //+ 
    18'h17437: Data = 4'h2; //+ 
    18'h17438: Data = 4'h2; //+ 
    18'h17439: Data = 4'h2; //+ 
    18'h17440: Data = 4'h2; //+ 
    18'h17441: Data = 4'h2; //+ 
    18'h17442: Data = 4'h2; //+ 
    18'h17443: Data = 4'h2; //+ 
    18'h17444: Data = 4'h2; //+ 
    18'h17445: Data = 4'h2; //+ 
    18'h17446: Data = 4'h6; //[ 
    18'h17447: Data = 4'h6; //[ 
    18'h17448: Data = 4'h4; //> 
    18'h17449: Data = 4'h4; //> 
    18'h17450: Data = 4'h4; //> 
    18'h17451: Data = 4'h4; //> 
    18'h17452: Data = 4'h4; //> 
    18'h17453: Data = 4'h4; //> 
    18'h17454: Data = 4'h4; //> 
    18'h17455: Data = 4'h4; //> 
    18'h17456: Data = 4'h4; //> 
    18'h17457: Data = 4'h7; //] 
    18'h17458: Data = 4'h2; //+ 
    18'h17459: Data = 4'h4; //> 
    18'h17460: Data = 4'ha; //0 
    18'h17461: Data = 4'h4; //> 
    18'h17462: Data = 4'ha; //0 
    18'h17463: Data = 4'h4; //> 
    18'h17464: Data = 4'ha; //0 
    18'h17465: Data = 4'h4; //> 
    18'h17466: Data = 4'ha; //0 
    18'h17467: Data = 4'h4; //> 
    18'h17468: Data = 4'ha; //0 
    18'h17469: Data = 4'h4; //> 
    18'h17470: Data = 4'ha; //0 
    18'h17471: Data = 4'h4; //> 
    18'h17472: Data = 4'ha; //0 
    18'h17473: Data = 4'h4; //> 
    18'h17474: Data = 4'ha; //0 
    18'h17475: Data = 4'h4; //> 
    18'h17476: Data = 4'ha; //0 
    18'h17477: Data = 4'h5; //< 
    18'h17478: Data = 4'h5; //< 
    18'h17479: Data = 4'h5; //< 
    18'h17480: Data = 4'h5; //< 
    18'h17481: Data = 4'h5; //< 
    18'h17482: Data = 4'h5; //< 
    18'h17483: Data = 4'h5; //< 
    18'h17484: Data = 4'h5; //< 
    18'h17485: Data = 4'h5; //< 
    18'h17486: Data = 4'h6; //[ 
    18'h17487: Data = 4'h5; //< 
    18'h17488: Data = 4'h5; //< 
    18'h17489: Data = 4'h5; //< 
    18'h17490: Data = 4'h5; //< 
    18'h17491: Data = 4'h5; //< 
    18'h17492: Data = 4'h5; //< 
    18'h17493: Data = 4'h5; //< 
    18'h17494: Data = 4'h5; //< 
    18'h17495: Data = 4'h5; //< 
    18'h17496: Data = 4'h7; //] 
    18'h17497: Data = 4'h4; //> 
    18'h17498: Data = 4'h4; //> 
    18'h17499: Data = 4'h4; //> 
    18'h17500: Data = 4'h4; //> 
    18'h17501: Data = 4'h4; //> 
    18'h17502: Data = 4'h4; //> 
    18'h17503: Data = 4'h4; //> 
    18'h17504: Data = 4'h4; //> 
    18'h17505: Data = 4'h4; //> 
    18'h17506: Data = 4'h3; //- 
    18'h17507: Data = 4'h7; //] 
    18'h17508: Data = 4'h2; //+ 
    18'h17509: Data = 4'h6; //[ 
    18'h17510: Data = 4'h4; //> 
    18'h17511: Data = 4'h2; //+ 
    18'h17512: Data = 4'h4; //> 
    18'h17513: Data = 4'h4; //> 
    18'h17514: Data = 4'h4; //> 
    18'h17515: Data = 4'h4; //> 
    18'h17516: Data = 4'h4; //> 
    18'h17517: Data = 4'h4; //> 
    18'h17518: Data = 4'h4; //> 
    18'h17519: Data = 4'h4; //> 
    18'h17520: Data = 4'h7; //] 
    18'h17521: Data = 4'h5; //< 
    18'h17522: Data = 4'h5; //< 
    18'h17523: Data = 4'h5; //< 
    18'h17524: Data = 4'h5; //< 
    18'h17525: Data = 4'h5; //< 
    18'h17526: Data = 4'h5; //< 
    18'h17527: Data = 4'h5; //< 
    18'h17528: Data = 4'h5; //< 
    18'h17529: Data = 4'h5; //< 
    18'h17530: Data = 4'h6; //[ 
    18'h17531: Data = 4'h5; //< 
    18'h17532: Data = 4'h5; //< 
    18'h17533: Data = 4'h5; //< 
    18'h17534: Data = 4'h5; //< 
    18'h17535: Data = 4'h5; //< 
    18'h17536: Data = 4'h5; //< 
    18'h17537: Data = 4'h5; //< 
    18'h17538: Data = 4'h5; //< 
    18'h17539: Data = 4'h5; //< 
    18'h17540: Data = 4'h7; //] 
    18'h17541: Data = 4'h4; //> 
    18'h17542: Data = 4'h4; //> 
    18'h17543: Data = 4'h4; //> 
    18'h17544: Data = 4'h4; //> 
    18'h17545: Data = 4'h4; //> 
    18'h17546: Data = 4'h4; //> 
    18'h17547: Data = 4'h4; //> 
    18'h17548: Data = 4'h4; //> 
    18'h17549: Data = 4'h4; //> 
    18'h17550: Data = 4'h6; //[ 
    18'h17551: Data = 4'h4; //> 
    18'h17552: Data = 4'h3; //- 
    18'h17553: Data = 4'h4; //> 
    18'h17554: Data = 4'h4; //> 
    18'h17555: Data = 4'h4; //> 
    18'h17556: Data = 4'h4; //> 
    18'h17557: Data = 4'h6; //[ 
    18'h17558: Data = 4'h3; //- 
    18'h17559: Data = 4'h5; //< 
    18'h17560: Data = 4'h5; //< 
    18'h17561: Data = 4'h5; //< 
    18'h17562: Data = 4'h5; //< 
    18'h17563: Data = 4'h2; //+ 
    18'h17564: Data = 4'h4; //> 
    18'h17565: Data = 4'h4; //> 
    18'h17566: Data = 4'h4; //> 
    18'h17567: Data = 4'h4; //> 
    18'h17568: Data = 4'h7; //] 
    18'h17569: Data = 4'h5; //< 
    18'h17570: Data = 4'h5; //< 
    18'h17571: Data = 4'h5; //< 
    18'h17572: Data = 4'h5; //< 
    18'h17573: Data = 4'h6; //[ 
    18'h17574: Data = 4'h3; //- 
    18'h17575: Data = 4'h4; //> 
    18'h17576: Data = 4'h4; //> 
    18'h17577: Data = 4'h4; //> 
    18'h17578: Data = 4'h4; //> 
    18'h17579: Data = 4'h2; //+ 
    18'h17580: Data = 4'h5; //< 
    18'h17581: Data = 4'h5; //< 
    18'h17582: Data = 4'h5; //< 
    18'h17583: Data = 4'h5; //< 
    18'h17584: Data = 4'h5; //< 
    18'h17585: Data = 4'h6; //[ 
    18'h17586: Data = 4'h3; //- 
    18'h17587: Data = 4'h4; //> 
    18'h17588: Data = 4'h4; //> 
    18'h17589: Data = 4'h6; //[ 
    18'h17590: Data = 4'h3; //- 
    18'h17591: Data = 4'h5; //< 
    18'h17592: Data = 4'h5; //< 
    18'h17593: Data = 4'h2; //+ 
    18'h17594: Data = 4'h4; //> 
    18'h17595: Data = 4'h4; //> 
    18'h17596: Data = 4'h7; //] 
    18'h17597: Data = 4'h5; //< 
    18'h17598: Data = 4'h5; //< 
    18'h17599: Data = 4'h6; //[ 
    18'h17600: Data = 4'h3; //- 
    18'h17601: Data = 4'h4; //> 
    18'h17602: Data = 4'h4; //> 
    18'h17603: Data = 4'h2; //+ 
    18'h17604: Data = 4'h4; //> 
    18'h17605: Data = 4'h4; //> 
    18'h17606: Data = 4'h2; //+ 
    18'h17607: Data = 4'h5; //< 
    18'h17608: Data = 4'h5; //< 
    18'h17609: Data = 4'h5; //< 
    18'h17610: Data = 4'h5; //< 
    18'h17611: Data = 4'h7; //] 
    18'h17612: Data = 4'h2; //+ 
    18'h17613: Data = 4'h4; //> 
    18'h17614: Data = 4'h4; //> 
    18'h17615: Data = 4'h4; //> 
    18'h17616: Data = 4'h4; //> 
    18'h17617: Data = 4'h4; //> 
    18'h17618: Data = 4'h4; //> 
    18'h17619: Data = 4'h4; //> 
    18'h17620: Data = 4'h4; //> 
    18'h17621: Data = 4'h4; //> 
    18'h17622: Data = 4'h7; //] 
    18'h17623: Data = 4'h5; //< 
    18'h17624: Data = 4'h5; //< 
    18'h17625: Data = 4'h5; //< 
    18'h17626: Data = 4'h5; //< 
    18'h17627: Data = 4'h5; //< 
    18'h17628: Data = 4'h5; //< 
    18'h17629: Data = 4'h5; //< 
    18'h17630: Data = 4'h5; //< 
    18'h17631: Data = 4'h6; //[ 
    18'h17632: Data = 4'h5; //< 
    18'h17633: Data = 4'h5; //< 
    18'h17634: Data = 4'h5; //< 
    18'h17635: Data = 4'h5; //< 
    18'h17636: Data = 4'h5; //< 
    18'h17637: Data = 4'h5; //< 
    18'h17638: Data = 4'h5; //< 
    18'h17639: Data = 4'h5; //< 
    18'h17640: Data = 4'h5; //< 
    18'h17641: Data = 4'h7; //] 
    18'h17642: Data = 4'h7; //] 
    18'h17643: Data = 4'h4; //> 
    18'h17644: Data = 4'h4; //> 
    18'h17645: Data = 4'h4; //> 
    18'h17646: Data = 4'h4; //> 
    18'h17647: Data = 4'h4; //> 
    18'h17648: Data = 4'h4; //> 
    18'h17649: Data = 4'h4; //> 
    18'h17650: Data = 4'h4; //> 
    18'h17651: Data = 4'h4; //> 
    18'h17652: Data = 4'h6; //[ 
    18'h17653: Data = 4'h4; //> 
    18'h17654: Data = 4'h4; //> 
    18'h17655: Data = 4'h4; //> 
    18'h17656: Data = 4'h4; //> 
    18'h17657: Data = 4'h4; //> 
    18'h17658: Data = 4'h4; //> 
    18'h17659: Data = 4'h4; //> 
    18'h17660: Data = 4'h4; //> 
    18'h17661: Data = 4'h4; //> 
    18'h17662: Data = 4'h7; //] 
    18'h17663: Data = 4'h5; //< 
    18'h17664: Data = 4'h5; //< 
    18'h17665: Data = 4'h5; //< 
    18'h17666: Data = 4'h5; //< 
    18'h17667: Data = 4'h5; //< 
    18'h17668: Data = 4'h5; //< 
    18'h17669: Data = 4'h5; //< 
    18'h17670: Data = 4'h5; //< 
    18'h17671: Data = 4'h5; //< 
    18'h17672: Data = 4'h6; //[ 
    18'h17673: Data = 4'h4; //> 
    18'h17674: Data = 4'h6; //[ 
    18'h17675: Data = 4'h3; //- 
    18'h17676: Data = 4'h4; //> 
    18'h17677: Data = 4'h4; //> 
    18'h17678: Data = 4'h4; //> 
    18'h17679: Data = 4'h4; //> 
    18'h17680: Data = 4'h4; //> 
    18'h17681: Data = 4'h4; //> 
    18'h17682: Data = 4'h4; //> 
    18'h17683: Data = 4'h4; //> 
    18'h17684: Data = 4'h4; //> 
    18'h17685: Data = 4'h2; //+ 
    18'h17686: Data = 4'h5; //< 
    18'h17687: Data = 4'h5; //< 
    18'h17688: Data = 4'h5; //< 
    18'h17689: Data = 4'h5; //< 
    18'h17690: Data = 4'h5; //< 
    18'h17691: Data = 4'h5; //< 
    18'h17692: Data = 4'h5; //< 
    18'h17693: Data = 4'h5; //< 
    18'h17694: Data = 4'h5; //< 
    18'h17695: Data = 4'h7; //] 
    18'h17696: Data = 4'h5; //< 
    18'h17697: Data = 4'h5; //< 
    18'h17698: Data = 4'h5; //< 
    18'h17699: Data = 4'h5; //< 
    18'h17700: Data = 4'h5; //< 
    18'h17701: Data = 4'h5; //< 
    18'h17702: Data = 4'h5; //< 
    18'h17703: Data = 4'h5; //< 
    18'h17704: Data = 4'h5; //< 
    18'h17705: Data = 4'h5; //< 
    18'h17706: Data = 4'h7; //] 
    18'h17707: Data = 4'h4; //> 
    18'h17708: Data = 4'h6; //[ 
    18'h17709: Data = 4'h3; //- 
    18'h17710: Data = 4'h4; //> 
    18'h17711: Data = 4'h4; //> 
    18'h17712: Data = 4'h4; //> 
    18'h17713: Data = 4'h4; //> 
    18'h17714: Data = 4'h4; //> 
    18'h17715: Data = 4'h4; //> 
    18'h17716: Data = 4'h4; //> 
    18'h17717: Data = 4'h4; //> 
    18'h17718: Data = 4'h4; //> 
    18'h17719: Data = 4'h2; //+ 
    18'h17720: Data = 4'h5; //< 
    18'h17721: Data = 4'h5; //< 
    18'h17722: Data = 4'h5; //< 
    18'h17723: Data = 4'h5; //< 
    18'h17724: Data = 4'h5; //< 
    18'h17725: Data = 4'h5; //< 
    18'h17726: Data = 4'h5; //< 
    18'h17727: Data = 4'h5; //< 
    18'h17728: Data = 4'h5; //< 
    18'h17729: Data = 4'h7; //] 
    18'h17730: Data = 4'h5; //< 
    18'h17731: Data = 4'h2; //+ 
    18'h17732: Data = 4'h4; //> 
    18'h17733: Data = 4'h4; //> 
    18'h17734: Data = 4'h4; //> 
    18'h17735: Data = 4'h4; //> 
    18'h17736: Data = 4'h4; //> 
    18'h17737: Data = 4'h4; //> 
    18'h17738: Data = 4'h4; //> 
    18'h17739: Data = 4'h4; //> 
    18'h17740: Data = 4'h7; //] 
    18'h17741: Data = 4'h5; //< 
    18'h17742: Data = 4'h5; //< 
    18'h17743: Data = 4'h5; //< 
    18'h17744: Data = 4'h5; //< 
    18'h17745: Data = 4'h5; //< 
    18'h17746: Data = 4'h5; //< 
    18'h17747: Data = 4'h5; //< 
    18'h17748: Data = 4'h5; //< 
    18'h17749: Data = 4'h5; //< 
    18'h17750: Data = 4'h6; //[ 
    18'h17751: Data = 4'h4; //> 
    18'h17752: Data = 4'h6; //[ 
    18'h17753: Data = 4'h3; //- 
    18'h17754: Data = 4'h7; //] 
    18'h17755: Data = 4'h5; //< 
    18'h17756: Data = 4'h3; //- 
    18'h17757: Data = 4'h4; //> 
    18'h17758: Data = 4'h4; //> 
    18'h17759: Data = 4'h4; //> 
    18'h17760: Data = 4'h4; //> 
    18'h17761: Data = 4'h6; //[ 
    18'h17762: Data = 4'h3; //- 
    18'h17763: Data = 4'h5; //< 
    18'h17764: Data = 4'h5; //< 
    18'h17765: Data = 4'h5; //< 
    18'h17766: Data = 4'h5; //< 
    18'h17767: Data = 4'h2; //+ 
    18'h17768: Data = 4'h4; //> 
    18'h17769: Data = 4'h6; //[ 
    18'h17770: Data = 4'h5; //< 
    18'h17771: Data = 4'h3; //- 
    18'h17772: Data = 4'h4; //> 
    18'h17773: Data = 4'h3; //- 
    18'h17774: Data = 4'h5; //< 
    18'h17775: Data = 4'h5; //< 
    18'h17776: Data = 4'h5; //< 
    18'h17777: Data = 4'h5; //< 
    18'h17778: Data = 4'h5; //< 
    18'h17779: Data = 4'h5; //< 
    18'h17780: Data = 4'h2; //+ 
    18'h17781: Data = 4'h4; //> 
    18'h17782: Data = 4'h4; //> 
    18'h17783: Data = 4'h4; //> 
    18'h17784: Data = 4'h4; //> 
    18'h17785: Data = 4'h4; //> 
    18'h17786: Data = 4'h4; //> 
    18'h17787: Data = 4'h7; //] 
    18'h17788: Data = 4'h5; //< 
    18'h17789: Data = 4'h6; //[ 
    18'h17790: Data = 4'h3; //- 
    18'h17791: Data = 4'h4; //> 
    18'h17792: Data = 4'h2; //+ 
    18'h17793: Data = 4'h5; //< 
    18'h17794: Data = 4'h7; //] 
    18'h17795: Data = 4'h4; //> 
    18'h17796: Data = 4'h4; //> 
    18'h17797: Data = 4'h4; //> 
    18'h17798: Data = 4'h4; //> 
    18'h17799: Data = 4'h7; //] 
    18'h17800: Data = 4'h5; //< 
    18'h17801: Data = 4'h5; //< 
    18'h17802: Data = 4'h5; //< 
    18'h17803: Data = 4'h6; //[ 
    18'h17804: Data = 4'h3; //- 
    18'h17805: Data = 4'h4; //> 
    18'h17806: Data = 4'h4; //> 
    18'h17807: Data = 4'h4; //> 
    18'h17808: Data = 4'h2; //+ 
    18'h17809: Data = 4'h5; //< 
    18'h17810: Data = 4'h5; //< 
    18'h17811: Data = 4'h5; //< 
    18'h17812: Data = 4'h7; //] 
    18'h17813: Data = 4'h5; //< 
    18'h17814: Data = 4'h2; //+ 
    18'h17815: Data = 4'h5; //< 
    18'h17816: Data = 4'h5; //< 
    18'h17817: Data = 4'h5; //< 
    18'h17818: Data = 4'h5; //< 
    18'h17819: Data = 4'h5; //< 
    18'h17820: Data = 4'h5; //< 
    18'h17821: Data = 4'h5; //< 
    18'h17822: Data = 4'h5; //< 
    18'h17823: Data = 4'h5; //< 
    18'h17824: Data = 4'h7; //] 
    18'h17825: Data = 4'h4; //> 
    18'h17826: Data = 4'h4; //> 
    18'h17827: Data = 4'h4; //> 
    18'h17828: Data = 4'h4; //> 
    18'h17829: Data = 4'h4; //> 
    18'h17830: Data = 4'h4; //> 
    18'h17831: Data = 4'h4; //> 
    18'h17832: Data = 4'h4; //> 
    18'h17833: Data = 4'h4; //> 
    18'h17834: Data = 4'h6; //[ 
    18'h17835: Data = 4'h4; //> 
    18'h17836: Data = 4'h2; //+ 
    18'h17837: Data = 4'h4; //> 
    18'h17838: Data = 4'h4; //> 
    18'h17839: Data = 4'h4; //> 
    18'h17840: Data = 4'h4; //> 
    18'h17841: Data = 4'h4; //> 
    18'h17842: Data = 4'h4; //> 
    18'h17843: Data = 4'h4; //> 
    18'h17844: Data = 4'h4; //> 
    18'h17845: Data = 4'h7; //] 
    18'h17846: Data = 4'h5; //< 
    18'h17847: Data = 4'h5; //< 
    18'h17848: Data = 4'h5; //< 
    18'h17849: Data = 4'h5; //< 
    18'h17850: Data = 4'h5; //< 
    18'h17851: Data = 4'h5; //< 
    18'h17852: Data = 4'h5; //< 
    18'h17853: Data = 4'h5; //< 
    18'h17854: Data = 4'h5; //< 
    18'h17855: Data = 4'h6; //[ 
    18'h17856: Data = 4'h5; //< 
    18'h17857: Data = 4'h5; //< 
    18'h17858: Data = 4'h5; //< 
    18'h17859: Data = 4'h5; //< 
    18'h17860: Data = 4'h5; //< 
    18'h17861: Data = 4'h5; //< 
    18'h17862: Data = 4'h5; //< 
    18'h17863: Data = 4'h5; //< 
    18'h17864: Data = 4'h5; //< 
    18'h17865: Data = 4'h7; //] 
    18'h17866: Data = 4'h4; //> 
    18'h17867: Data = 4'h4; //> 
    18'h17868: Data = 4'h4; //> 
    18'h17869: Data = 4'h4; //> 
    18'h17870: Data = 4'h4; //> 
    18'h17871: Data = 4'h4; //> 
    18'h17872: Data = 4'h4; //> 
    18'h17873: Data = 4'h4; //> 
    18'h17874: Data = 4'h4; //> 
    18'h17875: Data = 4'h6; //[ 
    18'h17876: Data = 4'h4; //> 
    18'h17877: Data = 4'h3; //- 
    18'h17878: Data = 4'h4; //> 
    18'h17879: Data = 4'h4; //> 
    18'h17880: Data = 4'h4; //> 
    18'h17881: Data = 4'h4; //> 
    18'h17882: Data = 4'h4; //> 
    18'h17883: Data = 4'h6; //[ 
    18'h17884: Data = 4'h3; //- 
    18'h17885: Data = 4'h5; //< 
    18'h17886: Data = 4'h5; //< 
    18'h17887: Data = 4'h5; //< 
    18'h17888: Data = 4'h5; //< 
    18'h17889: Data = 4'h5; //< 
    18'h17890: Data = 4'h2; //+ 
    18'h17891: Data = 4'h4; //> 
    18'h17892: Data = 4'h4; //> 
    18'h17893: Data = 4'h4; //> 
    18'h17894: Data = 4'h4; //> 
    18'h17895: Data = 4'h4; //> 
    18'h17896: Data = 4'h7; //] 
    18'h17897: Data = 4'h5; //< 
    18'h17898: Data = 4'h5; //< 
    18'h17899: Data = 4'h5; //< 
    18'h17900: Data = 4'h5; //< 
    18'h17901: Data = 4'h5; //< 
    18'h17902: Data = 4'h6; //[ 
    18'h17903: Data = 4'h3; //- 
    18'h17904: Data = 4'h4; //> 
    18'h17905: Data = 4'h4; //> 
    18'h17906: Data = 4'h4; //> 
    18'h17907: Data = 4'h4; //> 
    18'h17908: Data = 4'h4; //> 
    18'h17909: Data = 4'h2; //+ 
    18'h17910: Data = 4'h5; //< 
    18'h17911: Data = 4'h5; //< 
    18'h17912: Data = 4'h5; //< 
    18'h17913: Data = 4'h5; //< 
    18'h17914: Data = 4'h5; //< 
    18'h17915: Data = 4'h5; //< 
    18'h17916: Data = 4'h6; //[ 
    18'h17917: Data = 4'h3; //- 
    18'h17918: Data = 4'h4; //> 
    18'h17919: Data = 4'h4; //> 
    18'h17920: Data = 4'h4; //> 
    18'h17921: Data = 4'h6; //[ 
    18'h17922: Data = 4'h3; //- 
    18'h17923: Data = 4'h5; //< 
    18'h17924: Data = 4'h5; //< 
    18'h17925: Data = 4'h5; //< 
    18'h17926: Data = 4'h2; //+ 
    18'h17927: Data = 4'h4; //> 
    18'h17928: Data = 4'h4; //> 
    18'h17929: Data = 4'h4; //> 
    18'h17930: Data = 4'h7; //] 
    18'h17931: Data = 4'h5; //< 
    18'h17932: Data = 4'h5; //< 
    18'h17933: Data = 4'h5; //< 
    18'h17934: Data = 4'h6; //[ 
    18'h17935: Data = 4'h3; //- 
    18'h17936: Data = 4'h4; //> 
    18'h17937: Data = 4'h4; //> 
    18'h17938: Data = 4'h4; //> 
    18'h17939: Data = 4'h2; //+ 
    18'h17940: Data = 4'h4; //> 
    18'h17941: Data = 4'h2; //+ 
    18'h17942: Data = 4'h5; //< 
    18'h17943: Data = 4'h5; //< 
    18'h17944: Data = 4'h5; //< 
    18'h17945: Data = 4'h5; //< 
    18'h17946: Data = 4'h7; //] 
    18'h17947: Data = 4'h2; //+ 
    18'h17948: Data = 4'h4; //> 
    18'h17949: Data = 4'h4; //> 
    18'h17950: Data = 4'h4; //> 
    18'h17951: Data = 4'h4; //> 
    18'h17952: Data = 4'h4; //> 
    18'h17953: Data = 4'h4; //> 
    18'h17954: Data = 4'h4; //> 
    18'h17955: Data = 4'h4; //> 
    18'h17956: Data = 4'h4; //> 
    18'h17957: Data = 4'h7; //] 
    18'h17958: Data = 4'h5; //< 
    18'h17959: Data = 4'h5; //< 
    18'h17960: Data = 4'h5; //< 
    18'h17961: Data = 4'h5; //< 
    18'h17962: Data = 4'h5; //< 
    18'h17963: Data = 4'h5; //< 
    18'h17964: Data = 4'h5; //< 
    18'h17965: Data = 4'h5; //< 
    18'h17966: Data = 4'h6; //[ 
    18'h17967: Data = 4'h5; //< 
    18'h17968: Data = 4'h5; //< 
    18'h17969: Data = 4'h5; //< 
    18'h17970: Data = 4'h5; //< 
    18'h17971: Data = 4'h5; //< 
    18'h17972: Data = 4'h5; //< 
    18'h17973: Data = 4'h5; //< 
    18'h17974: Data = 4'h5; //< 
    18'h17975: Data = 4'h5; //< 
    18'h17976: Data = 4'h7; //] 
    18'h17977: Data = 4'h7; //] 
    18'h17978: Data = 4'h4; //> 
    18'h17979: Data = 4'h4; //> 
    18'h17980: Data = 4'h4; //> 
    18'h17981: Data = 4'h4; //> 
    18'h17982: Data = 4'h4; //> 
    18'h17983: Data = 4'h4; //> 
    18'h17984: Data = 4'h4; //> 
    18'h17985: Data = 4'h4; //> 
    18'h17986: Data = 4'h4; //> 
    18'h17987: Data = 4'h6; //[ 
    18'h17988: Data = 4'h4; //> 
    18'h17989: Data = 4'h4; //> 
    18'h17990: Data = 4'h4; //> 
    18'h17991: Data = 4'h4; //> 
    18'h17992: Data = 4'h4; //> 
    18'h17993: Data = 4'h4; //> 
    18'h17994: Data = 4'h4; //> 
    18'h17995: Data = 4'h4; //> 
    18'h17996: Data = 4'h4; //> 
    18'h17997: Data = 4'h7; //] 
    18'h17998: Data = 4'h5; //< 
    18'h17999: Data = 4'h5; //< 
    18'h18000: Data = 4'h5; //< 
    18'h18001: Data = 4'h5; //< 
    18'h18002: Data = 4'h5; //< 
    18'h18003: Data = 4'h5; //< 
    18'h18004: Data = 4'h5; //< 
    18'h18005: Data = 4'h5; //< 
    18'h18006: Data = 4'h5; //< 
    18'h18007: Data = 4'h6; //[ 
    18'h18008: Data = 4'h4; //> 
    18'h18009: Data = 4'h4; //> 
    18'h18010: Data = 4'h6; //[ 
    18'h18011: Data = 4'h3; //- 
    18'h18012: Data = 4'h4; //> 
    18'h18013: Data = 4'h4; //> 
    18'h18014: Data = 4'h4; //> 
    18'h18015: Data = 4'h4; //> 
    18'h18016: Data = 4'h4; //> 
    18'h18017: Data = 4'h4; //> 
    18'h18018: Data = 4'h4; //> 
    18'h18019: Data = 4'h4; //> 
    18'h18020: Data = 4'h4; //> 
    18'h18021: Data = 4'h2; //+ 
    18'h18022: Data = 4'h5; //< 
    18'h18023: Data = 4'h5; //< 
    18'h18024: Data = 4'h5; //< 
    18'h18025: Data = 4'h5; //< 
    18'h18026: Data = 4'h5; //< 
    18'h18027: Data = 4'h5; //< 
    18'h18028: Data = 4'h5; //< 
    18'h18029: Data = 4'h5; //< 
    18'h18030: Data = 4'h5; //< 
    18'h18031: Data = 4'h7; //] 
    18'h18032: Data = 4'h5; //< 
    18'h18033: Data = 4'h5; //< 
    18'h18034: Data = 4'h5; //< 
    18'h18035: Data = 4'h5; //< 
    18'h18036: Data = 4'h5; //< 
    18'h18037: Data = 4'h5; //< 
    18'h18038: Data = 4'h5; //< 
    18'h18039: Data = 4'h5; //< 
    18'h18040: Data = 4'h5; //< 
    18'h18041: Data = 4'h5; //< 
    18'h18042: Data = 4'h5; //< 
    18'h18043: Data = 4'h7; //] 
    18'h18044: Data = 4'h4; //> 
    18'h18045: Data = 4'h4; //> 
    18'h18046: Data = 4'h6; //[ 
    18'h18047: Data = 4'h3; //- 
    18'h18048: Data = 4'h4; //> 
    18'h18049: Data = 4'h4; //> 
    18'h18050: Data = 4'h4; //> 
    18'h18051: Data = 4'h4; //> 
    18'h18052: Data = 4'h4; //> 
    18'h18053: Data = 4'h4; //> 
    18'h18054: Data = 4'h4; //> 
    18'h18055: Data = 4'h4; //> 
    18'h18056: Data = 4'h4; //> 
    18'h18057: Data = 4'h2; //+ 
    18'h18058: Data = 4'h5; //< 
    18'h18059: Data = 4'h5; //< 
    18'h18060: Data = 4'h5; //< 
    18'h18061: Data = 4'h5; //< 
    18'h18062: Data = 4'h5; //< 
    18'h18063: Data = 4'h5; //< 
    18'h18064: Data = 4'h5; //< 
    18'h18065: Data = 4'h5; //< 
    18'h18066: Data = 4'h5; //< 
    18'h18067: Data = 4'h7; //] 
    18'h18068: Data = 4'h5; //< 
    18'h18069: Data = 4'h5; //< 
    18'h18070: Data = 4'h2; //+ 
    18'h18071: Data = 4'h4; //> 
    18'h18072: Data = 4'h4; //> 
    18'h18073: Data = 4'h4; //> 
    18'h18074: Data = 4'h4; //> 
    18'h18075: Data = 4'h4; //> 
    18'h18076: Data = 4'h4; //> 
    18'h18077: Data = 4'h4; //> 
    18'h18078: Data = 4'h4; //> 
    18'h18079: Data = 4'h7; //] 
    18'h18080: Data = 4'h5; //< 
    18'h18081: Data = 4'h5; //< 
    18'h18082: Data = 4'h5; //< 
    18'h18083: Data = 4'h5; //< 
    18'h18084: Data = 4'h5; //< 
    18'h18085: Data = 4'h5; //< 
    18'h18086: Data = 4'h5; //< 
    18'h18087: Data = 4'h5; //< 
    18'h18088: Data = 4'h5; //< 
    18'h18089: Data = 4'h6; //[ 
    18'h18090: Data = 4'h4; //> 
    18'h18091: Data = 4'ha; //0 
    18'h18092: Data = 4'h5; //< 
    18'h18093: Data = 4'h3; //- 
    18'h18094: Data = 4'h4; //> 
    18'h18095: Data = 4'h4; //> 
    18'h18096: Data = 4'h4; //> 
    18'h18097: Data = 4'h4; //> 
    18'h18098: Data = 4'h6; //[ 
    18'h18099: Data = 4'h3; //- 
    18'h18100: Data = 4'h5; //< 
    18'h18101: Data = 4'h5; //< 
    18'h18102: Data = 4'h5; //< 
    18'h18103: Data = 4'h5; //< 
    18'h18104: Data = 4'h2; //+ 
    18'h18105: Data = 4'h4; //> 
    18'h18106: Data = 4'h6; //[ 
    18'h18107: Data = 4'h5; //< 
    18'h18108: Data = 4'h3; //- 
    18'h18109: Data = 4'h4; //> 
    18'h18110: Data = 4'h3; //- 
    18'h18111: Data = 4'h5; //< 
    18'h18112: Data = 4'h5; //< 
    18'h18113: Data = 4'h5; //< 
    18'h18114: Data = 4'h5; //< 
    18'h18115: Data = 4'h5; //< 
    18'h18116: Data = 4'h5; //< 
    18'h18117: Data = 4'h2; //+ 
    18'h18118: Data = 4'h4; //> 
    18'h18119: Data = 4'h4; //> 
    18'h18120: Data = 4'h4; //> 
    18'h18121: Data = 4'h4; //> 
    18'h18122: Data = 4'h4; //> 
    18'h18123: Data = 4'h4; //> 
    18'h18124: Data = 4'h7; //] 
    18'h18125: Data = 4'h5; //< 
    18'h18126: Data = 4'h6; //[ 
    18'h18127: Data = 4'h3; //- 
    18'h18128: Data = 4'h4; //> 
    18'h18129: Data = 4'h2; //+ 
    18'h18130: Data = 4'h5; //< 
    18'h18131: Data = 4'h7; //] 
    18'h18132: Data = 4'h4; //> 
    18'h18133: Data = 4'h4; //> 
    18'h18134: Data = 4'h4; //> 
    18'h18135: Data = 4'h4; //> 
    18'h18136: Data = 4'h7; //] 
    18'h18137: Data = 4'h5; //< 
    18'h18138: Data = 4'h5; //< 
    18'h18139: Data = 4'h5; //< 
    18'h18140: Data = 4'h6; //[ 
    18'h18141: Data = 4'h3; //- 
    18'h18142: Data = 4'h4; //> 
    18'h18143: Data = 4'h4; //> 
    18'h18144: Data = 4'h4; //> 
    18'h18145: Data = 4'h2; //+ 
    18'h18146: Data = 4'h5; //< 
    18'h18147: Data = 4'h5; //< 
    18'h18148: Data = 4'h5; //< 
    18'h18149: Data = 4'h7; //] 
    18'h18150: Data = 4'h5; //< 
    18'h18151: Data = 4'h2; //+ 
    18'h18152: Data = 4'h5; //< 
    18'h18153: Data = 4'h5; //< 
    18'h18154: Data = 4'h5; //< 
    18'h18155: Data = 4'h5; //< 
    18'h18156: Data = 4'h5; //< 
    18'h18157: Data = 4'h5; //< 
    18'h18158: Data = 4'h5; //< 
    18'h18159: Data = 4'h5; //< 
    18'h18160: Data = 4'h5; //< 
    18'h18161: Data = 4'h7; //] 
    18'h18162: Data = 4'h4; //> 
    18'h18163: Data = 4'h4; //> 
    18'h18164: Data = 4'h4; //> 
    18'h18165: Data = 4'h4; //> 
    18'h18166: Data = 4'h4; //> 
    18'h18167: Data = 4'h4; //> 
    18'h18168: Data = 4'h4; //> 
    18'h18169: Data = 4'h4; //> 
    18'h18170: Data = 4'h4; //> 
    18'h18171: Data = 4'h6; //[ 
    18'h18172: Data = 4'h4; //> 
    18'h18173: Data = 4'h4; //> 
    18'h18174: Data = 4'h4; //> 
    18'h18175: Data = 4'h4; //> 
    18'h18176: Data = 4'h6; //[ 
    18'h18177: Data = 4'h3; //- 
    18'h18178: Data = 4'h5; //< 
    18'h18179: Data = 4'h5; //< 
    18'h18180: Data = 4'h5; //< 
    18'h18181: Data = 4'h5; //< 
    18'h18182: Data = 4'h5; //< 
    18'h18183: Data = 4'h5; //< 
    18'h18184: Data = 4'h5; //< 
    18'h18185: Data = 4'h5; //< 
    18'h18186: Data = 4'h5; //< 
    18'h18187: Data = 4'h5; //< 
    18'h18188: Data = 4'h5; //< 
    18'h18189: Data = 4'h5; //< 
    18'h18190: Data = 4'h5; //< 
    18'h18191: Data = 4'h5; //< 
    18'h18192: Data = 4'h5; //< 
    18'h18193: Data = 4'h5; //< 
    18'h18194: Data = 4'h5; //< 
    18'h18195: Data = 4'h5; //< 
    18'h18196: Data = 4'h5; //< 
    18'h18197: Data = 4'h5; //< 
    18'h18198: Data = 4'h5; //< 
    18'h18199: Data = 4'h5; //< 
    18'h18200: Data = 4'h5; //< 
    18'h18201: Data = 4'h5; //< 
    18'h18202: Data = 4'h5; //< 
    18'h18203: Data = 4'h5; //< 
    18'h18204: Data = 4'h5; //< 
    18'h18205: Data = 4'h5; //< 
    18'h18206: Data = 4'h5; //< 
    18'h18207: Data = 4'h5; //< 
    18'h18208: Data = 4'h5; //< 
    18'h18209: Data = 4'h5; //< 
    18'h18210: Data = 4'h5; //< 
    18'h18211: Data = 4'h5; //< 
    18'h18212: Data = 4'h5; //< 
    18'h18213: Data = 4'h5; //< 
    18'h18214: Data = 4'h2; //+ 
    18'h18215: Data = 4'h4; //> 
    18'h18216: Data = 4'h4; //> 
    18'h18217: Data = 4'h4; //> 
    18'h18218: Data = 4'h4; //> 
    18'h18219: Data = 4'h4; //> 
    18'h18220: Data = 4'h4; //> 
    18'h18221: Data = 4'h4; //> 
    18'h18222: Data = 4'h4; //> 
    18'h18223: Data = 4'h4; //> 
    18'h18224: Data = 4'h4; //> 
    18'h18225: Data = 4'h4; //> 
    18'h18226: Data = 4'h4; //> 
    18'h18227: Data = 4'h4; //> 
    18'h18228: Data = 4'h4; //> 
    18'h18229: Data = 4'h4; //> 
    18'h18230: Data = 4'h4; //> 
    18'h18231: Data = 4'h4; //> 
    18'h18232: Data = 4'h4; //> 
    18'h18233: Data = 4'h4; //> 
    18'h18234: Data = 4'h4; //> 
    18'h18235: Data = 4'h4; //> 
    18'h18236: Data = 4'h4; //> 
    18'h18237: Data = 4'h4; //> 
    18'h18238: Data = 4'h4; //> 
    18'h18239: Data = 4'h4; //> 
    18'h18240: Data = 4'h4; //> 
    18'h18241: Data = 4'h4; //> 
    18'h18242: Data = 4'h4; //> 
    18'h18243: Data = 4'h4; //> 
    18'h18244: Data = 4'h4; //> 
    18'h18245: Data = 4'h4; //> 
    18'h18246: Data = 4'h4; //> 
    18'h18247: Data = 4'h4; //> 
    18'h18248: Data = 4'h4; //> 
    18'h18249: Data = 4'h4; //> 
    18'h18250: Data = 4'h4; //> 
    18'h18251: Data = 4'h7; //] 
    18'h18252: Data = 4'h4; //> 
    18'h18253: Data = 4'h4; //> 
    18'h18254: Data = 4'h4; //> 
    18'h18255: Data = 4'h4; //> 
    18'h18256: Data = 4'h4; //> 
    18'h18257: Data = 4'h7; //] 
    18'h18258: Data = 4'h5; //< 
    18'h18259: Data = 4'h5; //< 
    18'h18260: Data = 4'h5; //< 
    18'h18261: Data = 4'h5; //< 
    18'h18262: Data = 4'h5; //< 
    18'h18263: Data = 4'h5; //< 
    18'h18264: Data = 4'h5; //< 
    18'h18265: Data = 4'h5; //< 
    18'h18266: Data = 4'h5; //< 
    18'h18267: Data = 4'h6; //[ 
    18'h18268: Data = 4'h5; //< 
    18'h18269: Data = 4'h5; //< 
    18'h18270: Data = 4'h5; //< 
    18'h18271: Data = 4'h5; //< 
    18'h18272: Data = 4'h5; //< 
    18'h18273: Data = 4'h5; //< 
    18'h18274: Data = 4'h5; //< 
    18'h18275: Data = 4'h5; //< 
    18'h18276: Data = 4'h5; //< 
    18'h18277: Data = 4'h7; //] 
    18'h18278: Data = 4'h4; //> 
    18'h18279: Data = 4'h4; //> 
    18'h18280: Data = 4'h4; //> 
    18'h18281: Data = 4'h4; //> 
    18'h18282: Data = 4'h4; //> 
    18'h18283: Data = 4'h4; //> 
    18'h18284: Data = 4'h4; //> 
    18'h18285: Data = 4'h4; //> 
    18'h18286: Data = 4'h4; //> 
    18'h18287: Data = 4'h2; //+ 
    18'h18288: Data = 4'h2; //+ 
    18'h18289: Data = 4'h2; //+ 
    18'h18290: Data = 4'h2; //+ 
    18'h18291: Data = 4'h2; //+ 
    18'h18292: Data = 4'h2; //+ 
    18'h18293: Data = 4'h2; //+ 
    18'h18294: Data = 4'h2; //+ 
    18'h18295: Data = 4'h2; //+ 
    18'h18296: Data = 4'h2; //+ 
    18'h18297: Data = 4'h2; //+ 
    18'h18298: Data = 4'h2; //+ 
    18'h18299: Data = 4'h2; //+ 
    18'h18300: Data = 4'h2; //+ 
    18'h18301: Data = 4'h2; //+ 
    18'h18302: Data = 4'h6; //[ 
    18'h18303: Data = 4'h6; //[ 
    18'h18304: Data = 4'h4; //> 
    18'h18305: Data = 4'h4; //> 
    18'h18306: Data = 4'h4; //> 
    18'h18307: Data = 4'h4; //> 
    18'h18308: Data = 4'h4; //> 
    18'h18309: Data = 4'h4; //> 
    18'h18310: Data = 4'h4; //> 
    18'h18311: Data = 4'h4; //> 
    18'h18312: Data = 4'h4; //> 
    18'h18313: Data = 4'h7; //] 
    18'h18314: Data = 4'h5; //< 
    18'h18315: Data = 4'h5; //< 
    18'h18316: Data = 4'h5; //< 
    18'h18317: Data = 4'h5; //< 
    18'h18318: Data = 4'h5; //< 
    18'h18319: Data = 4'h5; //< 
    18'h18320: Data = 4'h5; //< 
    18'h18321: Data = 4'h5; //< 
    18'h18322: Data = 4'h5; //< 
    18'h18323: Data = 4'h3; //- 
    18'h18324: Data = 4'h5; //< 
    18'h18325: Data = 4'h5; //< 
    18'h18326: Data = 4'h5; //< 
    18'h18327: Data = 4'h5; //< 
    18'h18328: Data = 4'h5; //< 
    18'h18329: Data = 4'h5; //< 
    18'h18330: Data = 4'h5; //< 
    18'h18331: Data = 4'h5; //< 
    18'h18332: Data = 4'h5; //< 
    18'h18333: Data = 4'h6; //[ 
    18'h18334: Data = 4'h5; //< 
    18'h18335: Data = 4'h5; //< 
    18'h18336: Data = 4'h5; //< 
    18'h18337: Data = 4'h5; //< 
    18'h18338: Data = 4'h5; //< 
    18'h18339: Data = 4'h5; //< 
    18'h18340: Data = 4'h5; //< 
    18'h18341: Data = 4'h5; //< 
    18'h18342: Data = 4'h5; //< 
    18'h18343: Data = 4'h7; //] 
    18'h18344: Data = 4'h4; //> 
    18'h18345: Data = 4'h4; //> 
    18'h18346: Data = 4'h4; //> 
    18'h18347: Data = 4'h4; //> 
    18'h18348: Data = 4'h4; //> 
    18'h18349: Data = 4'h4; //> 
    18'h18350: Data = 4'h4; //> 
    18'h18351: Data = 4'h4; //> 
    18'h18352: Data = 4'h4; //> 
    18'h18353: Data = 4'h3; //- 
    18'h18354: Data = 4'h7; //] 
    18'h18355: Data = 4'h2; //+ 
    18'h18356: Data = 4'h4; //> 
    18'h18357: Data = 4'h4; //> 
    18'h18358: Data = 4'h4; //> 
    18'h18359: Data = 4'h4; //> 
    18'h18360: Data = 4'h4; //> 
    18'h18361: Data = 4'h4; //> 
    18'h18362: Data = 4'h4; //> 
    18'h18363: Data = 4'h4; //> 
    18'h18364: Data = 4'h4; //> 
    18'h18365: Data = 4'h4; //> 
    18'h18366: Data = 4'h4; //> 
    18'h18367: Data = 4'h4; //> 
    18'h18368: Data = 4'h4; //> 
    18'h18369: Data = 4'h4; //> 
    18'h18370: Data = 4'h4; //> 
    18'h18371: Data = 4'h4; //> 
    18'h18372: Data = 4'h4; //> 
    18'h18373: Data = 4'h4; //> 
    18'h18374: Data = 4'h4; //> 
    18'h18375: Data = 4'h4; //> 
    18'h18376: Data = 4'h4; //> 
    18'h18377: Data = 4'h2; //+ 
    18'h18378: Data = 4'h5; //< 
    18'h18379: Data = 4'h5; //< 
    18'h18380: Data = 4'h5; //< 
    18'h18381: Data = 4'h6; //[ 
    18'h18382: Data = 4'h5; //< 
    18'h18383: Data = 4'h5; //< 
    18'h18384: Data = 4'h5; //< 
    18'h18385: Data = 4'h5; //< 
    18'h18386: Data = 4'h5; //< 
    18'h18387: Data = 4'h5; //< 
    18'h18388: Data = 4'h5; //< 
    18'h18389: Data = 4'h5; //< 
    18'h18390: Data = 4'h5; //< 
    18'h18391: Data = 4'h7; //] 
    18'h18392: Data = 4'h4; //> 
    18'h18393: Data = 4'h4; //> 
    18'h18394: Data = 4'h4; //> 
    18'h18395: Data = 4'h4; //> 
    18'h18396: Data = 4'h4; //> 
    18'h18397: Data = 4'h4; //> 
    18'h18398: Data = 4'h4; //> 
    18'h18399: Data = 4'h4; //> 
    18'h18400: Data = 4'h4; //> 
    18'h18401: Data = 4'h6; //[ 
    18'h18402: Data = 4'h4; //> 
    18'h18403: Data = 4'h4; //> 
    18'h18404: Data = 4'h4; //> 
    18'h18405: Data = 4'h6; //[ 
    18'h18406: Data = 4'h3; //- 
    18'h18407: Data = 4'h5; //< 
    18'h18408: Data = 4'h5; //< 
    18'h18409: Data = 4'h5; //< 
    18'h18410: Data = 4'h3; //- 
    18'h18411: Data = 4'h4; //> 
    18'h18412: Data = 4'h4; //> 
    18'h18413: Data = 4'h4; //> 
    18'h18414: Data = 4'h7; //] 
    18'h18415: Data = 4'h2; //+ 
    18'h18416: Data = 4'h5; //< 
    18'h18417: Data = 4'h5; //< 
    18'h18418: Data = 4'h5; //< 
    18'h18419: Data = 4'h6; //[ 
    18'h18420: Data = 4'h3; //- 
    18'h18421: Data = 4'h4; //> 
    18'h18422: Data = 4'h4; //> 
    18'h18423: Data = 4'h4; //> 
    18'h18424: Data = 4'h3; //- 
    18'h18425: Data = 4'h4; //> 
    18'h18426: Data = 4'h6; //[ 
    18'h18427: Data = 4'h3; //- 
    18'h18428: Data = 4'h5; //< 
    18'h18429: Data = 4'h5; //< 
    18'h18430: Data = 4'h5; //< 
    18'h18431: Data = 4'h5; //< 
    18'h18432: Data = 4'h2; //+ 
    18'h18433: Data = 4'h4; //> 
    18'h18434: Data = 4'h4; //> 
    18'h18435: Data = 4'h4; //> 
    18'h18436: Data = 4'h4; //> 
    18'h18437: Data = 4'h7; //] 
    18'h18438: Data = 4'h5; //< 
    18'h18439: Data = 4'h5; //< 
    18'h18440: Data = 4'h5; //< 
    18'h18441: Data = 4'h5; //< 
    18'h18442: Data = 4'h6; //[ 
    18'h18443: Data = 4'h3; //- 
    18'h18444: Data = 4'h4; //> 
    18'h18445: Data = 4'h4; //> 
    18'h18446: Data = 4'h4; //> 
    18'h18447: Data = 4'h4; //> 
    18'h18448: Data = 4'h2; //+ 
    18'h18449: Data = 4'h5; //< 
    18'h18450: Data = 4'h5; //< 
    18'h18451: Data = 4'h5; //< 
    18'h18452: Data = 4'h5; //< 
    18'h18453: Data = 4'h5; //< 
    18'h18454: Data = 4'h5; //< 
    18'h18455: Data = 4'h5; //< 
    18'h18456: Data = 4'h5; //< 
    18'h18457: Data = 4'h5; //< 
    18'h18458: Data = 4'h5; //< 
    18'h18459: Data = 4'h5; //< 
    18'h18460: Data = 4'h5; //< 
    18'h18461: Data = 4'h5; //< 
    18'h18462: Data = 4'h6; //[ 
    18'h18463: Data = 4'h5; //< 
    18'h18464: Data = 4'h5; //< 
    18'h18465: Data = 4'h5; //< 
    18'h18466: Data = 4'h5; //< 
    18'h18467: Data = 4'h5; //< 
    18'h18468: Data = 4'h5; //< 
    18'h18469: Data = 4'h5; //< 
    18'h18470: Data = 4'h5; //< 
    18'h18471: Data = 4'h5; //< 
    18'h18472: Data = 4'h7; //] 
    18'h18473: Data = 4'h4; //> 
    18'h18474: Data = 4'h4; //> 
    18'h18475: Data = 4'h4; //> 
    18'h18476: Data = 4'h4; //> 
    18'h18477: Data = 4'ha; //0 
    18'h18478: Data = 4'h2; //+ 
    18'h18479: Data = 4'h4; //> 
    18'h18480: Data = 4'h4; //> 
    18'h18481: Data = 4'h4; //> 
    18'h18482: Data = 4'h4; //> 
    18'h18483: Data = 4'h4; //> 
    18'h18484: Data = 4'h6; //[ 
    18'h18485: Data = 4'h4; //> 
    18'h18486: Data = 4'h4; //> 
    18'h18487: Data = 4'h4; //> 
    18'h18488: Data = 4'h4; //> 
    18'h18489: Data = 4'h4; //> 
    18'h18490: Data = 4'h4; //> 
    18'h18491: Data = 4'h4; //> 
    18'h18492: Data = 4'h4; //> 
    18'h18493: Data = 4'h4; //> 
    18'h18494: Data = 4'h7; //] 
    18'h18495: Data = 4'h4; //> 
    18'h18496: Data = 4'h2; //+ 
    18'h18497: Data = 4'h5; //< 
    18'h18498: Data = 4'h7; //] 
    18'h18499: Data = 4'h7; //] 
    18'h18500: Data = 4'h2; //+ 
    18'h18501: Data = 4'h4; //> 
    18'h18502: Data = 4'h4; //> 
    18'h18503: Data = 4'h4; //> 
    18'h18504: Data = 4'h4; //> 
    18'h18505: Data = 4'h6; //[ 
    18'h18506: Data = 4'h3; //- 
    18'h18507: Data = 4'h5; //< 
    18'h18508: Data = 4'h5; //< 
    18'h18509: Data = 4'h5; //< 
    18'h18510: Data = 4'h5; //< 
    18'h18511: Data = 4'h3; //- 
    18'h18512: Data = 4'h4; //> 
    18'h18513: Data = 4'h4; //> 
    18'h18514: Data = 4'h4; //> 
    18'h18515: Data = 4'h4; //> 
    18'h18516: Data = 4'h7; //] 
    18'h18517: Data = 4'h2; //+ 
    18'h18518: Data = 4'h5; //< 
    18'h18519: Data = 4'h5; //< 
    18'h18520: Data = 4'h5; //< 
    18'h18521: Data = 4'h5; //< 
    18'h18522: Data = 4'h6; //[ 
    18'h18523: Data = 4'h3; //- 
    18'h18524: Data = 4'h4; //> 
    18'h18525: Data = 4'h4; //> 
    18'h18526: Data = 4'h4; //> 
    18'h18527: Data = 4'h4; //> 
    18'h18528: Data = 4'h3; //- 
    18'h18529: Data = 4'h5; //< 
    18'h18530: Data = 4'h6; //[ 
    18'h18531: Data = 4'h3; //- 
    18'h18532: Data = 4'h5; //< 
    18'h18533: Data = 4'h5; //< 
    18'h18534: Data = 4'h5; //< 
    18'h18535: Data = 4'h2; //+ 
    18'h18536: Data = 4'h4; //> 
    18'h18537: Data = 4'h4; //> 
    18'h18538: Data = 4'h4; //> 
    18'h18539: Data = 4'h7; //] 
    18'h18540: Data = 4'h5; //< 
    18'h18541: Data = 4'h5; //< 
    18'h18542: Data = 4'h5; //< 
    18'h18543: Data = 4'h6; //[ 
    18'h18544: Data = 4'h3; //- 
    18'h18545: Data = 4'h4; //> 
    18'h18546: Data = 4'h4; //> 
    18'h18547: Data = 4'h4; //> 
    18'h18548: Data = 4'h2; //+ 
    18'h18549: Data = 4'h5; //< 
    18'h18550: Data = 4'h5; //< 
    18'h18551: Data = 4'h5; //< 
    18'h18552: Data = 4'h5; //< 
    18'h18553: Data = 4'h5; //< 
    18'h18554: Data = 4'h5; //< 
    18'h18555: Data = 4'h5; //< 
    18'h18556: Data = 4'h5; //< 
    18'h18557: Data = 4'h5; //< 
    18'h18558: Data = 4'h5; //< 
    18'h18559: Data = 4'h5; //< 
    18'h18560: Data = 4'h5; //< 
    18'h18561: Data = 4'h6; //[ 
    18'h18562: Data = 4'h5; //< 
    18'h18563: Data = 4'h5; //< 
    18'h18564: Data = 4'h5; //< 
    18'h18565: Data = 4'h5; //< 
    18'h18566: Data = 4'h5; //< 
    18'h18567: Data = 4'h5; //< 
    18'h18568: Data = 4'h5; //< 
    18'h18569: Data = 4'h5; //< 
    18'h18570: Data = 4'h5; //< 
    18'h18571: Data = 4'h7; //] 
    18'h18572: Data = 4'h4; //> 
    18'h18573: Data = 4'h4; //> 
    18'h18574: Data = 4'h4; //> 
    18'h18575: Data = 4'ha; //0 
    18'h18576: Data = 4'h2; //+ 
    18'h18577: Data = 4'h4; //> 
    18'h18578: Data = 4'h4; //> 
    18'h18579: Data = 4'h4; //> 
    18'h18580: Data = 4'h4; //> 
    18'h18581: Data = 4'h4; //> 
    18'h18582: Data = 4'h4; //> 
    18'h18583: Data = 4'h6; //[ 
    18'h18584: Data = 4'h4; //> 
    18'h18585: Data = 4'h4; //> 
    18'h18586: Data = 4'h4; //> 
    18'h18587: Data = 4'h4; //> 
    18'h18588: Data = 4'h4; //> 
    18'h18589: Data = 4'h4; //> 
    18'h18590: Data = 4'h4; //> 
    18'h18591: Data = 4'h4; //> 
    18'h18592: Data = 4'h4; //> 
    18'h18593: Data = 4'h7; //] 
    18'h18594: Data = 4'h4; //> 
    18'h18595: Data = 4'ha; //0 
    18'h18596: Data = 4'h2; //+ 
    18'h18597: Data = 4'h5; //< 
    18'h18598: Data = 4'h7; //] 
    18'h18599: Data = 4'h7; //] 
    18'h18600: Data = 4'h2; //+ 
    18'h18601: Data = 4'h4; //> 
    18'h18602: Data = 4'h6; //[ 
    18'h18603: Data = 4'h3; //- 
    18'h18604: Data = 4'h5; //< 
    18'h18605: Data = 4'h6; //[ 
    18'h18606: Data = 4'h4; //> 
    18'h18607: Data = 4'h4; //> 
    18'h18608: Data = 4'h4; //> 
    18'h18609: Data = 4'h4; //> 
    18'h18610: Data = 4'h4; //> 
    18'h18611: Data = 4'h4; //> 
    18'h18612: Data = 4'h4; //> 
    18'h18613: Data = 4'h4; //> 
    18'h18614: Data = 4'h4; //> 
    18'h18615: Data = 4'h7; //] 
    18'h18616: Data = 4'h5; //< 
    18'h18617: Data = 4'h5; //< 
    18'h18618: Data = 4'h5; //< 
    18'h18619: Data = 4'h5; //< 
    18'h18620: Data = 4'h5; //< 
    18'h18621: Data = 4'h5; //< 
    18'h18622: Data = 4'h5; //< 
    18'h18623: Data = 4'h5; //< 
    18'h18624: Data = 4'h7; //] 
    18'h18625: Data = 4'h4; //> 
    18'h18626: Data = 4'h4; //> 
    18'h18627: Data = 4'h4; //> 
    18'h18628: Data = 4'h4; //> 
    18'h18629: Data = 4'h4; //> 
    18'h18630: Data = 4'h4; //> 
    18'h18631: Data = 4'h4; //> 
    18'h18632: Data = 4'h4; //> 
    18'h18633: Data = 4'h7; //] 
    18'h18634: Data = 4'h5; //< 
    18'h18635: Data = 4'h5; //< 
    18'h18636: Data = 4'h5; //< 
    18'h18637: Data = 4'h5; //< 
    18'h18638: Data = 4'h5; //< 
    18'h18639: Data = 4'h5; //< 
    18'h18640: Data = 4'h5; //< 
    18'h18641: Data = 4'h5; //< 
    18'h18642: Data = 4'h5; //< 
    18'h18643: Data = 4'h6; //[ 
    18'h18644: Data = 4'h5; //< 
    18'h18645: Data = 4'h5; //< 
    18'h18646: Data = 4'h5; //< 
    18'h18647: Data = 4'h5; //< 
    18'h18648: Data = 4'h5; //< 
    18'h18649: Data = 4'h5; //< 
    18'h18650: Data = 4'h5; //< 
    18'h18651: Data = 4'h5; //< 
    18'h18652: Data = 4'h5; //< 
    18'h18653: Data = 4'h7; //] 
    18'h18654: Data = 4'h4; //> 
    18'h18655: Data = 4'h4; //> 
    18'h18656: Data = 4'h3; //- 
    18'h18657: Data = 4'h4; //> 
    18'h18658: Data = 4'h4; //> 
    18'h18659: Data = 4'h6; //[ 
    18'h18660: Data = 4'h3; //- 
    18'h18661: Data = 4'h5; //< 
    18'h18662: Data = 4'h5; //< 
    18'h18663: Data = 4'h5; //< 
    18'h18664: Data = 4'h5; //< 
    18'h18665: Data = 4'h2; //+ 
    18'h18666: Data = 4'h4; //> 
    18'h18667: Data = 4'h4; //> 
    18'h18668: Data = 4'h4; //> 
    18'h18669: Data = 4'h4; //> 
    18'h18670: Data = 4'h7; //] 
    18'h18671: Data = 4'h5; //< 
    18'h18672: Data = 4'h5; //< 
    18'h18673: Data = 4'h5; //< 
    18'h18674: Data = 4'h5; //< 
    18'h18675: Data = 4'h6; //[ 
    18'h18676: Data = 4'h3; //- 
    18'h18677: Data = 4'h4; //> 
    18'h18678: Data = 4'h4; //> 
    18'h18679: Data = 4'h4; //> 
    18'h18680: Data = 4'h4; //> 
    18'h18681: Data = 4'h2; //+ 
    18'h18682: Data = 4'h5; //< 
    18'h18683: Data = 4'h5; //< 
    18'h18684: Data = 4'ha; //0 
    18'h18685: Data = 4'h5; //< 
    18'h18686: Data = 4'h5; //< 
    18'h18687: Data = 4'h7; //] 
    18'h18688: Data = 4'h4; //> 
    18'h18689: Data = 4'h4; //> 
    18'h18690: Data = 4'h7; //] 
    18'h18691: Data = 4'h5; //< 
    18'h18692: Data = 4'h5; //< 
    18'h18693: Data = 4'h2; //+ 
    18'h18694: Data = 4'h4; //> 
    18'h18695: Data = 4'h4; //> 
    18'h18696: Data = 4'h4; //> 
    18'h18697: Data = 4'h4; //> 
    18'h18698: Data = 4'h6; //[ 
    18'h18699: Data = 4'h3; //- 
    18'h18700: Data = 4'h5; //< 
    18'h18701: Data = 4'h5; //< 
    18'h18702: Data = 4'h5; //< 
    18'h18703: Data = 4'h5; //< 
    18'h18704: Data = 4'h3; //- 
    18'h18705: Data = 4'h4; //> 
    18'h18706: Data = 4'h4; //> 
    18'h18707: Data = 4'h4; //> 
    18'h18708: Data = 4'h4; //> 
    18'h18709: Data = 4'h7; //] 
    18'h18710: Data = 4'h2; //+ 
    18'h18711: Data = 4'h5; //< 
    18'h18712: Data = 4'h5; //< 
    18'h18713: Data = 4'h5; //< 
    18'h18714: Data = 4'h5; //< 
    18'h18715: Data = 4'h6; //[ 
    18'h18716: Data = 4'h3; //- 
    18'h18717: Data = 4'h4; //> 
    18'h18718: Data = 4'h4; //> 
    18'h18719: Data = 4'h4; //> 
    18'h18720: Data = 4'h4; //> 
    18'h18721: Data = 4'h3; //- 
    18'h18722: Data = 4'h5; //< 
    18'h18723: Data = 4'h5; //< 
    18'h18724: Data = 4'h5; //< 
    18'h18725: Data = 4'h5; //< 
    18'h18726: Data = 4'h5; //< 
    18'h18727: Data = 4'h5; //< 
    18'h18728: Data = 4'h8; //. 
    18'h18729: Data = 4'h4; //> 
    18'h18730: Data = 4'h4; //> 
    18'h18731: Data = 4'h7; //] 
    18'h18732: Data = 4'h4; //> 
    18'h18733: Data = 4'h4; //> 
    18'h18734: Data = 4'h4; //> 
    18'h18735: Data = 4'h4; //> 
    18'h18736: Data = 4'h6; //[ 
    18'h18737: Data = 4'h3; //- 
    18'h18738: Data = 4'h5; //< 
    18'h18739: Data = 4'h5; //< 
    18'h18740: Data = 4'h5; //< 
    18'h18741: Data = 4'h5; //< 
    18'h18742: Data = 4'h5; //< 
    18'h18743: Data = 4'h5; //< 
    18'h18744: Data = 4'h5; //< 
    18'h18745: Data = 4'h8; //. 
    18'h18746: Data = 4'h4; //> 
    18'h18747: Data = 4'h4; //> 
    18'h18748: Data = 4'h4; //> 
    18'h18749: Data = 4'h4; //> 
    18'h18750: Data = 4'h4; //> 
    18'h18751: Data = 4'h4; //> 
    18'h18752: Data = 4'h4; //> 
    18'h18753: Data = 4'h7; //] 
    18'h18754: Data = 4'h5; //< 
    18'h18755: Data = 4'h5; //< 
    18'h18756: Data = 4'h5; //< 
    18'h18757: Data = 4'ha; //0 
    18'h18758: Data = 4'h4; //> 
    18'h18759: Data = 4'ha; //0 
    18'h18760: Data = 4'h4; //> 
    18'h18761: Data = 4'ha; //0 
    18'h18762: Data = 4'h4; //> 
    18'h18763: Data = 4'ha; //0 
    18'h18764: Data = 4'h4; //> 
    18'h18765: Data = 4'ha; //0 
    18'h18766: Data = 4'h4; //> 
    18'h18767: Data = 4'ha; //0 
    18'h18768: Data = 4'h4; //> 
    18'h18769: Data = 4'h4; //> 
    18'h18770: Data = 4'h4; //> 
    18'h18771: Data = 4'h6; //[ 
    18'h18772: Data = 4'h4; //> 
    18'h18773: Data = 4'ha; //0 
    18'h18774: Data = 4'h4; //> 
    18'h18775: Data = 4'ha; //0 
    18'h18776: Data = 4'h4; //> 
    18'h18777: Data = 4'ha; //0 
    18'h18778: Data = 4'h4; //> 
    18'h18779: Data = 4'ha; //0 
    18'h18780: Data = 4'h4; //> 
    18'h18781: Data = 4'ha; //0 
    18'h18782: Data = 4'h4; //> 
    18'h18783: Data = 4'ha; //0 
    18'h18784: Data = 4'h4; //> 
    18'h18785: Data = 4'h4; //> 
    18'h18786: Data = 4'h4; //> 
    18'h18787: Data = 4'h7; //] 
    18'h18788: Data = 4'h5; //< 
    18'h18789: Data = 4'h5; //< 
    18'h18790: Data = 4'h5; //< 
    18'h18791: Data = 4'h5; //< 
    18'h18792: Data = 4'h5; //< 
    18'h18793: Data = 4'h5; //< 
    18'h18794: Data = 4'h5; //< 
    18'h18795: Data = 4'h5; //< 
    18'h18796: Data = 4'h5; //< 
    18'h18797: Data = 4'h6; //[ 
    18'h18798: Data = 4'h5; //< 
    18'h18799: Data = 4'h5; //< 
    18'h18800: Data = 4'h5; //< 
    18'h18801: Data = 4'h5; //< 
    18'h18802: Data = 4'h5; //< 
    18'h18803: Data = 4'h5; //< 
    18'h18804: Data = 4'h5; //< 
    18'h18805: Data = 4'h5; //< 
    18'h18806: Data = 4'h5; //< 
    18'h18807: Data = 4'h7; //] 
    18'h18808: Data = 4'h4; //> 
    18'h18809: Data = 4'h4; //> 
    18'h18810: Data = 4'h4; //> 
    18'h18811: Data = 4'h4; //> 
    18'h18812: Data = 4'h4; //> 
    18'h18813: Data = 4'h4; //> 
    18'h18814: Data = 4'h4; //> 
    18'h18815: Data = 4'h4; //> 
    18'h18816: Data = 4'h4; //> 
    18'h18817: Data = 4'h6; //[ 
    18'h18818: Data = 4'h4; //> 
    18'h18819: Data = 4'h4; //> 
    18'h18820: Data = 4'h4; //> 
    18'h18821: Data = 4'h4; //> 
    18'h18822: Data = 4'h4; //> 
    18'h18823: Data = 4'ha; //0 
    18'h18824: Data = 4'h4; //> 
    18'h18825: Data = 4'h4; //> 
    18'h18826: Data = 4'h4; //> 
    18'h18827: Data = 4'h4; //> 
    18'h18828: Data = 4'h7; //] 
    18'h18829: Data = 4'h5; //< 
    18'h18830: Data = 4'h5; //< 
    18'h18831: Data = 4'h5; //< 
    18'h18832: Data = 4'h5; //< 
    18'h18833: Data = 4'h5; //< 
    18'h18834: Data = 4'h5; //< 
    18'h18835: Data = 4'h5; //< 
    18'h18836: Data = 4'h5; //< 
    18'h18837: Data = 4'h5; //< 
    18'h18838: Data = 4'h6; //[ 
    18'h18839: Data = 4'h5; //< 
    18'h18840: Data = 4'h5; //< 
    18'h18841: Data = 4'h5; //< 
    18'h18842: Data = 4'h5; //< 
    18'h18843: Data = 4'h5; //< 
    18'h18844: Data = 4'h5; //< 
    18'h18845: Data = 4'h5; //< 
    18'h18846: Data = 4'h5; //< 
    18'h18847: Data = 4'h5; //< 
    18'h18848: Data = 4'h7; //] 
    18'h18849: Data = 4'h4; //> 
    18'h18850: Data = 4'h2; //+ 
    18'h18851: Data = 4'h2; //+ 
    18'h18852: Data = 4'h2; //+ 
    18'h18853: Data = 4'h2; //+ 
    18'h18854: Data = 4'h2; //+ 
    18'h18855: Data = 4'h2; //+ 
    18'h18856: Data = 4'h2; //+ 
    18'h18857: Data = 4'h2; //+ 
    18'h18858: Data = 4'h2; //+ 
    18'h18859: Data = 4'h2; //+ 
    18'h18860: Data = 4'h2; //+ 
    18'h18861: Data = 4'h6; //[ 
    18'h18862: Data = 4'h3; //- 
    18'h18863: Data = 4'h6; //[ 
    18'h18864: Data = 4'h3; //- 
    18'h18865: Data = 4'h4; //> 
    18'h18866: Data = 4'h4; //> 
    18'h18867: Data = 4'h4; //> 
    18'h18868: Data = 4'h4; //> 
    18'h18869: Data = 4'h4; //> 
    18'h18870: Data = 4'h4; //> 
    18'h18871: Data = 4'h4; //> 
    18'h18872: Data = 4'h4; //> 
    18'h18873: Data = 4'h4; //> 
    18'h18874: Data = 4'h2; //+ 
    18'h18875: Data = 4'h5; //< 
    18'h18876: Data = 4'h5; //< 
    18'h18877: Data = 4'h5; //< 
    18'h18878: Data = 4'h5; //< 
    18'h18879: Data = 4'h5; //< 
    18'h18880: Data = 4'h5; //< 
    18'h18881: Data = 4'h5; //< 
    18'h18882: Data = 4'h5; //< 
    18'h18883: Data = 4'h5; //< 
    18'h18884: Data = 4'h7; //] 
    18'h18885: Data = 4'h4; //> 
    18'h18886: Data = 4'h4; //> 
    18'h18887: Data = 4'h4; //> 
    18'h18888: Data = 4'h4; //> 
    18'h18889: Data = 4'h4; //> 
    18'h18890: Data = 4'h4; //> 
    18'h18891: Data = 4'h4; //> 
    18'h18892: Data = 4'h4; //> 
    18'h18893: Data = 4'h4; //> 
    18'h18894: Data = 4'h7; //] 
    18'h18895: Data = 4'h4; //> 
    18'h18896: Data = 4'h4; //> 
    18'h18897: Data = 4'h4; //> 
    18'h18898: Data = 4'h4; //> 
    18'h18899: Data = 4'h2; //+ 
    18'h18900: Data = 4'h4; //> 
    18'h18901: Data = 4'h4; //> 
    18'h18902: Data = 4'h4; //> 
    18'h18903: Data = 4'h4; //> 
    18'h18904: Data = 4'h4; //> 
    18'h18905: Data = 4'h4; //> 
    18'h18906: Data = 4'h4; //> 
    18'h18907: Data = 4'h4; //> 
    18'h18908: Data = 4'h4; //> 
    18'h18909: Data = 4'h2; //+ 
    18'h18910: Data = 4'h5; //< 
    18'h18911: Data = 4'h5; //< 
    18'h18912: Data = 4'h5; //< 
    18'h18913: Data = 4'h5; //< 
    18'h18914: Data = 4'h5; //< 
    18'h18915: Data = 4'h5; //< 
    18'h18916: Data = 4'h5; //< 
    18'h18917: Data = 4'h5; //< 
    18'h18918: Data = 4'h5; //< 
    18'h18919: Data = 4'h5; //< 
    18'h18920: Data = 4'h5; //< 
    18'h18921: Data = 4'h5; //< 
    18'h18922: Data = 4'h5; //< 
    18'h18923: Data = 4'h5; //< 
    18'h18924: Data = 4'h6; //[ 
    18'h18925: Data = 4'h5; //< 
    18'h18926: Data = 4'h5; //< 
    18'h18927: Data = 4'h5; //< 
    18'h18928: Data = 4'h5; //< 
    18'h18929: Data = 4'h5; //< 
    18'h18930: Data = 4'h5; //< 
    18'h18931: Data = 4'h5; //< 
    18'h18932: Data = 4'h5; //< 
    18'h18933: Data = 4'h5; //< 
    18'h18934: Data = 4'h7; //] 
    18'h18935: Data = 4'h4; //> 
    18'h18936: Data = 4'h4; //> 
    18'h18937: Data = 4'h4; //> 
    18'h18938: Data = 4'h4; //> 
    18'h18939: Data = 4'h4; //> 
    18'h18940: Data = 4'h4; //> 
    18'h18941: Data = 4'h4; //> 
    18'h18942: Data = 4'h6; //[ 
    18'h18943: Data = 4'h3; //- 
    18'h18944: Data = 4'h5; //< 
    18'h18945: Data = 4'h5; //< 
    18'h18946: Data = 4'h5; //< 
    18'h18947: Data = 4'h5; //< 
    18'h18948: Data = 4'h5; //< 
    18'h18949: Data = 4'h5; //< 
    18'h18950: Data = 4'h5; //< 
    18'h18951: Data = 4'h2; //+ 
    18'h18952: Data = 4'h4; //> 
    18'h18953: Data = 4'h4; //> 
    18'h18954: Data = 4'h4; //> 
    18'h18955: Data = 4'h4; //> 
    18'h18956: Data = 4'h4; //> 
    18'h18957: Data = 4'h4; //> 
    18'h18958: Data = 4'h4; //> 
    18'h18959: Data = 4'h7; //] 
    18'h18960: Data = 4'h5; //< 
    18'h18961: Data = 4'h5; //< 
    18'h18962: Data = 4'h5; //< 
    18'h18963: Data = 4'h5; //< 
    18'h18964: Data = 4'h5; //< 
    18'h18965: Data = 4'h5; //< 
    18'h18966: Data = 4'h5; //< 
    18'h18967: Data = 4'h6; //[ 
    18'h18968: Data = 4'h3; //- 
    18'h18969: Data = 4'h4; //> 
    18'h18970: Data = 4'h4; //> 
    18'h18971: Data = 4'h4; //> 
    18'h18972: Data = 4'h4; //> 
    18'h18973: Data = 4'h4; //> 
    18'h18974: Data = 4'h4; //> 
    18'h18975: Data = 4'h4; //> 
    18'h18976: Data = 4'h2; //+ 
    18'h18977: Data = 4'ha; //0 
    18'h18978: Data = 4'h4; //> 
    18'h18979: Data = 4'h4; //> 
    18'h18980: Data = 4'h6; //[ 
    18'h18981: Data = 4'h4; //> 
    18'h18982: Data = 4'h4; //> 
    18'h18983: Data = 4'h4; //> 
    18'h18984: Data = 4'h4; //> 
    18'h18985: Data = 4'h4; //> 
    18'h18986: Data = 4'h4; //> 
    18'h18987: Data = 4'h4; //> 
    18'h18988: Data = 4'h4; //> 
    18'h18989: Data = 4'h4; //> 
    18'h18990: Data = 4'h7; //] 
    18'h18991: Data = 4'h5; //< 
    18'h18992: Data = 4'h5; //< 
    18'h18993: Data = 4'h5; //< 
    18'h18994: Data = 4'h5; //< 
    18'h18995: Data = 4'h5; //< 
    18'h18996: Data = 4'h5; //< 
    18'h18997: Data = 4'h5; //< 
    18'h18998: Data = 4'h5; //< 
    18'h18999: Data = 4'h5; //< 
    18'h19000: Data = 4'h6; //[ 
    18'h19001: Data = 4'h4; //> 
    18'h19002: Data = 4'h4; //> 
    18'h19003: Data = 4'h4; //> 
    18'h19004: Data = 4'h4; //> 
    18'h19005: Data = 4'h4; //> 
    18'h19006: Data = 4'h4; //> 
    18'h19007: Data = 4'h4; //> 
    18'h19008: Data = 4'h6; //[ 
    18'h19009: Data = 4'h3; //- 
    18'h19010: Data = 4'h5; //< 
    18'h19011: Data = 4'h5; //< 
    18'h19012: Data = 4'h5; //< 
    18'h19013: Data = 4'h5; //< 
    18'h19014: Data = 4'h5; //< 
    18'h19015: Data = 4'h5; //< 
    18'h19016: Data = 4'h2; //+ 
    18'h19017: Data = 4'h4; //> 
    18'h19018: Data = 4'h4; //> 
    18'h19019: Data = 4'h4; //> 
    18'h19020: Data = 4'h4; //> 
    18'h19021: Data = 4'h4; //> 
    18'h19022: Data = 4'h4; //> 
    18'h19023: Data = 4'h7; //] 
    18'h19024: Data = 4'h5; //< 
    18'h19025: Data = 4'h5; //< 
    18'h19026: Data = 4'h5; //< 
    18'h19027: Data = 4'h5; //< 
    18'h19028: Data = 4'h5; //< 
    18'h19029: Data = 4'h5; //< 
    18'h19030: Data = 4'h6; //[ 
    18'h19031: Data = 4'h3; //- 
    18'h19032: Data = 4'h4; //> 
    18'h19033: Data = 4'h4; //> 
    18'h19034: Data = 4'h4; //> 
    18'h19035: Data = 4'h4; //> 
    18'h19036: Data = 4'h4; //> 
    18'h19037: Data = 4'h4; //> 
    18'h19038: Data = 4'h2; //+ 
    18'h19039: Data = 4'h5; //< 
    18'h19040: Data = 4'h5; //< 
    18'h19041: Data = 4'h5; //< 
    18'h19042: Data = 4'h5; //< 
    18'h19043: Data = 4'h5; //< 
    18'h19044: Data = 4'h5; //< 
    18'h19045: Data = 4'h5; //< 
    18'h19046: Data = 4'h6; //[ 
    18'h19047: Data = 4'h5; //< 
    18'h19048: Data = 4'h5; //< 
    18'h19049: Data = 4'h5; //< 
    18'h19050: Data = 4'h5; //< 
    18'h19051: Data = 4'h5; //< 
    18'h19052: Data = 4'h5; //< 
    18'h19053: Data = 4'h5; //< 
    18'h19054: Data = 4'h5; //< 
    18'h19055: Data = 4'h5; //< 
    18'h19056: Data = 4'h7; //] 
    18'h19057: Data = 4'h4; //> 
    18'h19058: Data = 4'h4; //> 
    18'h19059: Data = 4'h4; //> 
    18'h19060: Data = 4'h4; //> 
    18'h19061: Data = 4'h4; //> 
    18'h19062: Data = 4'h4; //> 
    18'h19063: Data = 4'h4; //> 
    18'h19064: Data = 4'ha; //0 
    18'h19065: Data = 4'h2; //+ 
    18'h19066: Data = 4'h4; //> 
    18'h19067: Data = 4'h4; //> 
    18'h19068: Data = 4'h4; //> 
    18'h19069: Data = 4'h7; //] 
    18'h19070: Data = 4'h5; //< 
    18'h19071: Data = 4'h5; //< 
    18'h19072: Data = 4'h5; //< 
    18'h19073: Data = 4'h5; //< 
    18'h19074: Data = 4'h5; //< 
    18'h19075: Data = 4'h5; //< 
    18'h19076: Data = 4'h5; //< 
    18'h19077: Data = 4'h5; //< 
    18'h19078: Data = 4'h5; //< 
    18'h19079: Data = 4'h5; //< 
    18'h19080: Data = 4'h7; //] 
    18'h19081: Data = 4'h7; //] 
    18'h19082: Data = 4'h4; //> 
    18'h19083: Data = 4'h4; //> 
    18'h19084: Data = 4'h4; //> 
    18'h19085: Data = 4'h4; //> 
    18'h19086: Data = 4'h4; //> 
    18'h19087: Data = 4'h4; //> 
    18'h19088: Data = 4'h4; //> 
    18'h19089: Data = 4'h6; //[ 
    18'h19090: Data = 4'h3; //- 
    18'h19091: Data = 4'h5; //< 
    18'h19092: Data = 4'h5; //< 
    18'h19093: Data = 4'h5; //< 
    18'h19094: Data = 4'h5; //< 
    18'h19095: Data = 4'h5; //< 
    18'h19096: Data = 4'h5; //< 
    18'h19097: Data = 4'h5; //< 
    18'h19098: Data = 4'h2; //+ 
    18'h19099: Data = 4'h4; //> 
    18'h19100: Data = 4'h4; //> 
    18'h19101: Data = 4'h4; //> 
    18'h19102: Data = 4'h4; //> 
    18'h19103: Data = 4'h4; //> 
    18'h19104: Data = 4'h4; //> 
    18'h19105: Data = 4'h4; //> 
    18'h19106: Data = 4'h7; //] 
    18'h19107: Data = 4'h5; //< 
    18'h19108: Data = 4'h5; //< 
    18'h19109: Data = 4'h5; //< 
    18'h19110: Data = 4'h5; //< 
    18'h19111: Data = 4'h5; //< 
    18'h19112: Data = 4'h5; //< 
    18'h19113: Data = 4'h5; //< 
    18'h19114: Data = 4'h6; //[ 
    18'h19115: Data = 4'h3; //- 
    18'h19116: Data = 4'h4; //> 
    18'h19117: Data = 4'h4; //> 
    18'h19118: Data = 4'h4; //> 
    18'h19119: Data = 4'h4; //> 
    18'h19120: Data = 4'h4; //> 
    18'h19121: Data = 4'h4; //> 
    18'h19122: Data = 4'h4; //> 
    18'h19123: Data = 4'h2; //+ 
    18'h19124: Data = 4'h4; //> 
    18'h19125: Data = 4'h4; //> 
    18'h19126: Data = 4'h6; //[ 
    18'h19127: Data = 4'h4; //> 
    18'h19128: Data = 4'h2; //+ 
    18'h19129: Data = 4'h4; //> 
    18'h19130: Data = 4'h4; //> 
    18'h19131: Data = 4'h4; //> 
    18'h19132: Data = 4'h4; //> 
    18'h19133: Data = 4'h6; //[ 
    18'h19134: Data = 4'h3; //- 
    18'h19135: Data = 4'h5; //< 
    18'h19136: Data = 4'h5; //< 
    18'h19137: Data = 4'h5; //< 
    18'h19138: Data = 4'h5; //< 
    18'h19139: Data = 4'h3; //- 
    18'h19140: Data = 4'h4; //> 
    18'h19141: Data = 4'h4; //> 
    18'h19142: Data = 4'h4; //> 
    18'h19143: Data = 4'h4; //> 
    18'h19144: Data = 4'h7; //] 
    18'h19145: Data = 4'h5; //< 
    18'h19146: Data = 4'h5; //< 
    18'h19147: Data = 4'h5; //< 
    18'h19148: Data = 4'h5; //< 
    18'h19149: Data = 4'h6; //[ 
    18'h19150: Data = 4'h3; //- 
    18'h19151: Data = 4'h4; //> 
    18'h19152: Data = 4'h4; //> 
    18'h19153: Data = 4'h4; //> 
    18'h19154: Data = 4'h4; //> 
    18'h19155: Data = 4'h2; //+ 
    18'h19156: Data = 4'h5; //< 
    18'h19157: Data = 4'h5; //< 
    18'h19158: Data = 4'h5; //< 
    18'h19159: Data = 4'h5; //< 
    18'h19160: Data = 4'h7; //] 
    18'h19161: Data = 4'h4; //> 
    18'h19162: Data = 4'h4; //> 
    18'h19163: Data = 4'h4; //> 
    18'h19164: Data = 4'h4; //> 
    18'h19165: Data = 4'h4; //> 
    18'h19166: Data = 4'h4; //> 
    18'h19167: Data = 4'h4; //> 
    18'h19168: Data = 4'h4; //> 
    18'h19169: Data = 4'h7; //] 
    18'h19170: Data = 4'h5; //< 
    18'h19171: Data = 4'h5; //< 
    18'h19172: Data = 4'h2; //+ 
    18'h19173: Data = 4'h5; //< 
    18'h19174: Data = 4'h5; //< 
    18'h19175: Data = 4'h5; //< 
    18'h19176: Data = 4'h5; //< 
    18'h19177: Data = 4'h5; //< 
    18'h19178: Data = 4'h5; //< 
    18'h19179: Data = 4'h5; //< 
    18'h19180: Data = 4'h6; //[ 
    18'h19181: Data = 4'h4; //> 
    18'h19182: Data = 4'h4; //> 
    18'h19183: Data = 4'h4; //> 
    18'h19184: Data = 4'h4; //> 
    18'h19185: Data = 4'h4; //> 
    18'h19186: Data = 4'h6; //[ 
    18'h19187: Data = 4'h3; //- 
    18'h19188: Data = 4'h4; //> 
    18'h19189: Data = 4'h4; //> 
    18'h19190: Data = 4'h2; //+ 
    18'h19191: Data = 4'h5; //< 
    18'h19192: Data = 4'h5; //< 
    18'h19193: Data = 4'h7; //] 
    18'h19194: Data = 4'h5; //< 
    18'h19195: Data = 4'h5; //< 
    18'h19196: Data = 4'h5; //< 
    18'h19197: Data = 4'h5; //< 
    18'h19198: Data = 4'h5; //< 
    18'h19199: Data = 4'h5; //< 
    18'h19200: Data = 4'h5; //< 
    18'h19201: Data = 4'h5; //< 
    18'h19202: Data = 4'h5; //< 
    18'h19203: Data = 4'h5; //< 
    18'h19204: Data = 4'h5; //< 
    18'h19205: Data = 4'h5; //< 
    18'h19206: Data = 4'h5; //< 
    18'h19207: Data = 4'h5; //< 
    18'h19208: Data = 4'h7; //] 
    18'h19209: Data = 4'h4; //> 
    18'h19210: Data = 4'h4; //> 
    18'h19211: Data = 4'h4; //> 
    18'h19212: Data = 4'h4; //> 
    18'h19213: Data = 4'h4; //> 
    18'h19214: Data = 4'h4; //> 
    18'h19215: Data = 4'h4; //> 
    18'h19216: Data = 4'h4; //> 
    18'h19217: Data = 4'h4; //> 
    18'h19218: Data = 4'h6; //[ 
    18'h19219: Data = 4'h4; //> 
    18'h19220: Data = 4'h4; //> 
    18'h19221: Data = 4'h4; //> 
    18'h19222: Data = 4'h4; //> 
    18'h19223: Data = 4'h4; //> 
    18'h19224: Data = 4'h4; //> 
    18'h19225: Data = 4'h4; //> 
    18'h19226: Data = 4'h4; //> 
    18'h19227: Data = 4'h4; //> 
    18'h19228: Data = 4'h7; //] 
    18'h19229: Data = 4'h5; //< 
    18'h19230: Data = 4'h5; //< 
    18'h19231: Data = 4'h5; //< 
    18'h19232: Data = 4'h5; //< 
    18'h19233: Data = 4'h5; //< 
    18'h19234: Data = 4'h5; //< 
    18'h19235: Data = 4'h5; //< 
    18'h19236: Data = 4'h5; //< 
    18'h19237: Data = 4'h5; //< 
    18'h19238: Data = 4'h6; //[ 
    18'h19239: Data = 4'h4; //> 
    18'h19240: Data = 4'ha; //0 
    18'h19241: Data = 4'h5; //< 
    18'h19242: Data = 4'h3; //- 
    18'h19243: Data = 4'h4; //> 
    18'h19244: Data = 4'h4; //> 
    18'h19245: Data = 4'h4; //> 
    18'h19246: Data = 4'h4; //> 
    18'h19247: Data = 4'h4; //> 
    18'h19248: Data = 4'h4; //> 
    18'h19249: Data = 4'h4; //> 
    18'h19250: Data = 4'h6; //[ 
    18'h19251: Data = 4'h3; //- 
    18'h19252: Data = 4'h5; //< 
    18'h19253: Data = 4'h5; //< 
    18'h19254: Data = 4'h5; //< 
    18'h19255: Data = 4'h5; //< 
    18'h19256: Data = 4'h5; //< 
    18'h19257: Data = 4'h5; //< 
    18'h19258: Data = 4'h5; //< 
    18'h19259: Data = 4'h2; //+ 
    18'h19260: Data = 4'h4; //> 
    18'h19261: Data = 4'h6; //[ 
    18'h19262: Data = 4'h5; //< 
    18'h19263: Data = 4'h3; //- 
    18'h19264: Data = 4'h4; //> 
    18'h19265: Data = 4'h3; //- 
    18'h19266: Data = 4'h5; //< 
    18'h19267: Data = 4'h5; //< 
    18'h19268: Data = 4'h5; //< 
    18'h19269: Data = 4'h2; //+ 
    18'h19270: Data = 4'h4; //> 
    18'h19271: Data = 4'h4; //> 
    18'h19272: Data = 4'h4; //> 
    18'h19273: Data = 4'h7; //] 
    18'h19274: Data = 4'h5; //< 
    18'h19275: Data = 4'h6; //[ 
    18'h19276: Data = 4'h3; //- 
    18'h19277: Data = 4'h4; //> 
    18'h19278: Data = 4'h2; //+ 
    18'h19279: Data = 4'h5; //< 
    18'h19280: Data = 4'h7; //] 
    18'h19281: Data = 4'h4; //> 
    18'h19282: Data = 4'h4; //> 
    18'h19283: Data = 4'h4; //> 
    18'h19284: Data = 4'h4; //> 
    18'h19285: Data = 4'h4; //> 
    18'h19286: Data = 4'h4; //> 
    18'h19287: Data = 4'h4; //> 
    18'h19288: Data = 4'h7; //] 
    18'h19289: Data = 4'h5; //< 
    18'h19290: Data = 4'h5; //< 
    18'h19291: Data = 4'h5; //< 
    18'h19292: Data = 4'h5; //< 
    18'h19293: Data = 4'h5; //< 
    18'h19294: Data = 4'h5; //< 
    18'h19295: Data = 4'h6; //[ 
    18'h19296: Data = 4'h3; //- 
    18'h19297: Data = 4'h4; //> 
    18'h19298: Data = 4'h4; //> 
    18'h19299: Data = 4'h4; //> 
    18'h19300: Data = 4'h4; //> 
    18'h19301: Data = 4'h4; //> 
    18'h19302: Data = 4'h4; //> 
    18'h19303: Data = 4'h2; //+ 
    18'h19304: Data = 4'h5; //< 
    18'h19305: Data = 4'h5; //< 
    18'h19306: Data = 4'h5; //< 
    18'h19307: Data = 4'h5; //< 
    18'h19308: Data = 4'h5; //< 
    18'h19309: Data = 4'h5; //< 
    18'h19310: Data = 4'h7; //] 
    18'h19311: Data = 4'h5; //< 
    18'h19312: Data = 4'h2; //+ 
    18'h19313: Data = 4'h5; //< 
    18'h19314: Data = 4'h5; //< 
    18'h19315: Data = 4'h5; //< 
    18'h19316: Data = 4'h5; //< 
    18'h19317: Data = 4'h5; //< 
    18'h19318: Data = 4'h5; //< 
    18'h19319: Data = 4'h5; //< 
    18'h19320: Data = 4'h5; //< 
    18'h19321: Data = 4'h5; //< 
    18'h19322: Data = 4'h7; //] 
    18'h19323: Data = 4'h4; //> 
    18'h19324: Data = 4'h4; //> 
    18'h19325: Data = 4'h4; //> 
    18'h19326: Data = 4'h4; //> 
    18'h19327: Data = 4'h4; //> 
    18'h19328: Data = 4'h4; //> 
    18'h19329: Data = 4'h4; //> 
    18'h19330: Data = 4'h3; //- 
    18'h19331: Data = 4'h5; //< 
    18'h19332: Data = 4'h5; //< 
    18'h19333: Data = 4'h5; //< 
    18'h19334: Data = 4'h5; //< 
    18'h19335: Data = 4'ha; //0 
    18'h19336: Data = 4'h2; //+ 
    18'h19337: Data = 4'h5; //< 
    18'h19338: Data = 4'h5; //< 
    18'h19339: Data = 4'h5; //< 
    18'h19340: Data = 4'h7; //] 
    18'h19341: Data = 4'h2; //+ 
    18'h19342: Data = 4'h4; //> 
    18'h19343: Data = 4'h4; //> 
    18'h19344: Data = 4'h4; //> 
    18'h19345: Data = 4'h4; //> 
    18'h19346: Data = 4'h4; //> 
    18'h19347: Data = 4'h4; //> 
    18'h19348: Data = 4'h4; //> 
    18'h19349: Data = 4'h6; //[ 
    18'h19350: Data = 4'h3; //- 
    18'h19351: Data = 4'h5; //< 
    18'h19352: Data = 4'h5; //< 
    18'h19353: Data = 4'h5; //< 
    18'h19354: Data = 4'h5; //< 
    18'h19355: Data = 4'h5; //< 
    18'h19356: Data = 4'h5; //< 
    18'h19357: Data = 4'h5; //< 
    18'h19358: Data = 4'h3; //- 
    18'h19359: Data = 4'h4; //> 
    18'h19360: Data = 4'h4; //> 
    18'h19361: Data = 4'h4; //> 
    18'h19362: Data = 4'h4; //> 
    18'h19363: Data = 4'h4; //> 
    18'h19364: Data = 4'h4; //> 
    18'h19365: Data = 4'h4; //> 
    18'h19366: Data = 4'h7; //] 
    18'h19367: Data = 4'h2; //+ 
    18'h19368: Data = 4'h5; //< 
    18'h19369: Data = 4'h5; //< 
    18'h19370: Data = 4'h5; //< 
    18'h19371: Data = 4'h5; //< 
    18'h19372: Data = 4'h5; //< 
    18'h19373: Data = 4'h5; //< 
    18'h19374: Data = 4'h5; //< 
    18'h19375: Data = 4'h6; //[ 
    18'h19376: Data = 4'h3; //- 
    18'h19377: Data = 4'h4; //> 
    18'h19378: Data = 4'h4; //> 
    18'h19379: Data = 4'h4; //> 
    18'h19380: Data = 4'h4; //> 
    18'h19381: Data = 4'h4; //> 
    18'h19382: Data = 4'h4; //> 
    18'h19383: Data = 4'h4; //> 
    18'h19384: Data = 4'h3; //- 
    18'h19385: Data = 4'h4; //> 
    18'h19386: Data = 4'h4; //> 
    18'h19387: Data = 4'h6; //[ 
    18'h19388: Data = 4'h4; //> 
    18'h19389: Data = 4'h4; //> 
    18'h19390: Data = 4'h4; //> 
    18'h19391: Data = 4'h4; //> 
    18'h19392: Data = 4'h4; //> 
    18'h19393: Data = 4'h6; //[ 
    18'h19394: Data = 4'h3; //- 
    18'h19395: Data = 4'h4; //> 
    18'h19396: Data = 4'h4; //> 
    18'h19397: Data = 4'h2; //+ 
    18'h19398: Data = 4'h5; //< 
    18'h19399: Data = 4'h5; //< 
    18'h19400: Data = 4'h7; //] 
    18'h19401: Data = 4'h4; //> 
    18'h19402: Data = 4'h4; //> 
    18'h19403: Data = 4'h4; //> 
    18'h19404: Data = 4'h4; //> 
    18'h19405: Data = 4'h7; //] 
    18'h19406: Data = 4'h5; //< 
    18'h19407: Data = 4'h5; //< 
    18'h19408: Data = 4'h5; //< 
    18'h19409: Data = 4'h5; //< 
    18'h19410: Data = 4'h5; //< 
    18'h19411: Data = 4'h5; //< 
    18'h19412: Data = 4'h5; //< 
    18'h19413: Data = 4'h5; //< 
    18'h19414: Data = 4'h5; //< 
    18'h19415: Data = 4'h6; //[ 
    18'h19416: Data = 4'h4; //> 
    18'h19417: Data = 4'ha; //0 
    18'h19418: Data = 4'h5; //< 
    18'h19419: Data = 4'h3; //- 
    18'h19420: Data = 4'h4; //> 
    18'h19421: Data = 4'h4; //> 
    18'h19422: Data = 4'h4; //> 
    18'h19423: Data = 4'h4; //> 
    18'h19424: Data = 4'h4; //> 
    18'h19425: Data = 4'h4; //> 
    18'h19426: Data = 4'h4; //> 
    18'h19427: Data = 4'h6; //[ 
    18'h19428: Data = 4'h3; //- 
    18'h19429: Data = 4'h5; //< 
    18'h19430: Data = 4'h5; //< 
    18'h19431: Data = 4'h5; //< 
    18'h19432: Data = 4'h5; //< 
    18'h19433: Data = 4'h5; //< 
    18'h19434: Data = 4'h5; //< 
    18'h19435: Data = 4'h5; //< 
    18'h19436: Data = 4'h2; //+ 
    18'h19437: Data = 4'h4; //> 
    18'h19438: Data = 4'h6; //[ 
    18'h19439: Data = 4'h5; //< 
    18'h19440: Data = 4'h3; //- 
    18'h19441: Data = 4'h4; //> 
    18'h19442: Data = 4'h3; //- 
    18'h19443: Data = 4'h5; //< 
    18'h19444: Data = 4'h5; //< 
    18'h19445: Data = 4'h5; //< 
    18'h19446: Data = 4'h2; //+ 
    18'h19447: Data = 4'h4; //> 
    18'h19448: Data = 4'h4; //> 
    18'h19449: Data = 4'h4; //> 
    18'h19450: Data = 4'h7; //] 
    18'h19451: Data = 4'h5; //< 
    18'h19452: Data = 4'h6; //[ 
    18'h19453: Data = 4'h3; //- 
    18'h19454: Data = 4'h4; //> 
    18'h19455: Data = 4'h2; //+ 
    18'h19456: Data = 4'h5; //< 
    18'h19457: Data = 4'h7; //] 
    18'h19458: Data = 4'h4; //> 
    18'h19459: Data = 4'h4; //> 
    18'h19460: Data = 4'h4; //> 
    18'h19461: Data = 4'h4; //> 
    18'h19462: Data = 4'h4; //> 
    18'h19463: Data = 4'h4; //> 
    18'h19464: Data = 4'h4; //> 
    18'h19465: Data = 4'h7; //] 
    18'h19466: Data = 4'h5; //< 
    18'h19467: Data = 4'h5; //< 
    18'h19468: Data = 4'h5; //< 
    18'h19469: Data = 4'h5; //< 
    18'h19470: Data = 4'h5; //< 
    18'h19471: Data = 4'h5; //< 
    18'h19472: Data = 4'h6; //[ 
    18'h19473: Data = 4'h3; //- 
    18'h19474: Data = 4'h4; //> 
    18'h19475: Data = 4'h4; //> 
    18'h19476: Data = 4'h4; //> 
    18'h19477: Data = 4'h4; //> 
    18'h19478: Data = 4'h4; //> 
    18'h19479: Data = 4'h4; //> 
    18'h19480: Data = 4'h2; //+ 
    18'h19481: Data = 4'h5; //< 
    18'h19482: Data = 4'h5; //< 
    18'h19483: Data = 4'h5; //< 
    18'h19484: Data = 4'h5; //< 
    18'h19485: Data = 4'h5; //< 
    18'h19486: Data = 4'h5; //< 
    18'h19487: Data = 4'h7; //] 
    18'h19488: Data = 4'h5; //< 
    18'h19489: Data = 4'h2; //+ 
    18'h19490: Data = 4'h5; //< 
    18'h19491: Data = 4'h5; //< 
    18'h19492: Data = 4'h5; //< 
    18'h19493: Data = 4'h5; //< 
    18'h19494: Data = 4'h5; //< 
    18'h19495: Data = 4'h5; //< 
    18'h19496: Data = 4'h5; //< 
    18'h19497: Data = 4'h5; //< 
    18'h19498: Data = 4'h5; //< 
    18'h19499: Data = 4'h7; //] 
    18'h19500: Data = 4'h4; //> 
    18'h19501: Data = 4'h2; //+ 
    18'h19502: Data = 4'h2; //+ 
    18'h19503: Data = 4'h2; //+ 
    18'h19504: Data = 4'h2; //+ 
    18'h19505: Data = 4'h2; //+ 
    18'h19506: Data = 4'h6; //[ 
    18'h19507: Data = 4'h3; //- 
    18'h19508: Data = 4'h6; //[ 
    18'h19509: Data = 4'h3; //- 
    18'h19510: Data = 4'h4; //> 
    18'h19511: Data = 4'h4; //> 
    18'h19512: Data = 4'h4; //> 
    18'h19513: Data = 4'h4; //> 
    18'h19514: Data = 4'h4; //> 
    18'h19515: Data = 4'h4; //> 
    18'h19516: Data = 4'h4; //> 
    18'h19517: Data = 4'h4; //> 
    18'h19518: Data = 4'h4; //> 
    18'h19519: Data = 4'h2; //+ 
    18'h19520: Data = 4'h5; //< 
    18'h19521: Data = 4'h5; //< 
    18'h19522: Data = 4'h5; //< 
    18'h19523: Data = 4'h5; //< 
    18'h19524: Data = 4'h5; //< 
    18'h19525: Data = 4'h5; //< 
    18'h19526: Data = 4'h5; //< 
    18'h19527: Data = 4'h5; //< 
    18'h19528: Data = 4'h5; //< 
    18'h19529: Data = 4'h7; //] 
    18'h19530: Data = 4'h4; //> 
    18'h19531: Data = 4'h4; //> 
    18'h19532: Data = 4'h4; //> 
    18'h19533: Data = 4'h4; //> 
    18'h19534: Data = 4'h4; //> 
    18'h19535: Data = 4'h4; //> 
    18'h19536: Data = 4'h4; //> 
    18'h19537: Data = 4'h4; //> 
    18'h19538: Data = 4'h4; //> 
    18'h19539: Data = 4'h7; //] 
    18'h19540: Data = 4'h4; //> 
    18'h19541: Data = 4'h4; //> 
    18'h19542: Data = 4'h4; //> 
    18'h19543: Data = 4'h4; //> 
    18'h19544: Data = 4'h2; //+ 
    18'h19545: Data = 4'h5; //< 
    18'h19546: Data = 4'h5; //< 
    18'h19547: Data = 4'h5; //< 
    18'h19548: Data = 4'h5; //< 
    18'h19549: Data = 4'h5; //< 
    18'h19550: Data = 4'h6; //[ 
    18'h19551: Data = 4'h5; //< 
    18'h19552: Data = 4'h5; //< 
    18'h19553: Data = 4'h5; //< 
    18'h19554: Data = 4'h5; //< 
    18'h19555: Data = 4'h5; //< 
    18'h19556: Data = 4'h5; //< 
    18'h19557: Data = 4'h5; //< 
    18'h19558: Data = 4'h5; //< 
    18'h19559: Data = 4'h5; //< 
    18'h19560: Data = 4'h7; //] 
    18'h19561: Data = 4'h4; //> 
    18'h19562: Data = 4'h4; //> 
    18'h19563: Data = 4'h4; //> 
    18'h19564: Data = 4'h4; //> 
    18'h19565: Data = 4'h4; //> 
    18'h19566: Data = 4'h4; //> 
    18'h19567: Data = 4'h4; //> 
    18'h19568: Data = 4'h4; //> 
    18'h19569: Data = 4'h4; //> 
    18'h19570: Data = 4'h6; //[ 
    18'h19571: Data = 4'h4; //> 
    18'h19572: Data = 4'h4; //> 
    18'h19573: Data = 4'h4; //> 
    18'h19574: Data = 4'h4; //> 
    18'h19575: Data = 4'h4; //> 
    18'h19576: Data = 4'h6; //[ 
    18'h19577: Data = 4'h3; //- 
    18'h19578: Data = 4'h5; //< 
    18'h19579: Data = 4'h5; //< 
    18'h19580: Data = 4'h5; //< 
    18'h19581: Data = 4'h5; //< 
    18'h19582: Data = 4'h5; //< 
    18'h19583: Data = 4'h3; //- 
    18'h19584: Data = 4'h4; //> 
    18'h19585: Data = 4'h4; //> 
    18'h19586: Data = 4'h4; //> 
    18'h19587: Data = 4'h4; //> 
    18'h19588: Data = 4'h4; //> 
    18'h19589: Data = 4'h7; //] 
    18'h19590: Data = 4'h2; //+ 
    18'h19591: Data = 4'h5; //< 
    18'h19592: Data = 4'h5; //< 
    18'h19593: Data = 4'h5; //< 
    18'h19594: Data = 4'h5; //< 
    18'h19595: Data = 4'h5; //< 
    18'h19596: Data = 4'h6; //[ 
    18'h19597: Data = 4'h3; //- 
    18'h19598: Data = 4'h4; //> 
    18'h19599: Data = 4'h4; //> 
    18'h19600: Data = 4'h4; //> 
    18'h19601: Data = 4'h4; //> 
    18'h19602: Data = 4'h4; //> 
    18'h19603: Data = 4'h3; //- 
    18'h19604: Data = 4'h4; //> 
    18'h19605: Data = 4'h4; //> 
    18'h19606: Data = 4'h6; //[ 
    18'h19607: Data = 4'h3; //- 
    18'h19608: Data = 4'h5; //< 
    18'h19609: Data = 4'h5; //< 
    18'h19610: Data = 4'h5; //< 
    18'h19611: Data = 4'h5; //< 
    18'h19612: Data = 4'h5; //< 
    18'h19613: Data = 4'h5; //< 
    18'h19614: Data = 4'h5; //< 
    18'h19615: Data = 4'h2; //+ 
    18'h19616: Data = 4'h4; //> 
    18'h19617: Data = 4'h4; //> 
    18'h19618: Data = 4'h4; //> 
    18'h19619: Data = 4'h4; //> 
    18'h19620: Data = 4'h4; //> 
    18'h19621: Data = 4'h4; //> 
    18'h19622: Data = 4'h4; //> 
    18'h19623: Data = 4'h7; //] 
    18'h19624: Data = 4'h5; //< 
    18'h19625: Data = 4'h5; //< 
    18'h19626: Data = 4'h5; //< 
    18'h19627: Data = 4'h5; //< 
    18'h19628: Data = 4'h5; //< 
    18'h19629: Data = 4'h5; //< 
    18'h19630: Data = 4'h5; //< 
    18'h19631: Data = 4'h6; //[ 
    18'h19632: Data = 4'h3; //- 
    18'h19633: Data = 4'h4; //> 
    18'h19634: Data = 4'h4; //> 
    18'h19635: Data = 4'h4; //> 
    18'h19636: Data = 4'h4; //> 
    18'h19637: Data = 4'h4; //> 
    18'h19638: Data = 4'h4; //> 
    18'h19639: Data = 4'h4; //> 
    18'h19640: Data = 4'h2; //+ 
    18'h19641: Data = 4'h5; //< 
    18'h19642: Data = 4'h5; //< 
    18'h19643: Data = 4'h5; //< 
    18'h19644: Data = 4'h5; //< 
    18'h19645: Data = 4'h5; //< 
    18'h19646: Data = 4'h5; //< 
    18'h19647: Data = 4'h5; //< 
    18'h19648: Data = 4'h5; //< 
    18'h19649: Data = 4'h5; //< 
    18'h19650: Data = 4'h5; //< 
    18'h19651: Data = 4'h5; //< 
    18'h19652: Data = 4'h5; //< 
    18'h19653: Data = 4'h5; //< 
    18'h19654: Data = 4'h5; //< 
    18'h19655: Data = 4'h5; //< 
    18'h19656: Data = 4'h5; //< 
    18'h19657: Data = 4'h6; //[ 
    18'h19658: Data = 4'h5; //< 
    18'h19659: Data = 4'h5; //< 
    18'h19660: Data = 4'h5; //< 
    18'h19661: Data = 4'h5; //< 
    18'h19662: Data = 4'h5; //< 
    18'h19663: Data = 4'h5; //< 
    18'h19664: Data = 4'h5; //< 
    18'h19665: Data = 4'h5; //< 
    18'h19666: Data = 4'h5; //< 
    18'h19667: Data = 4'h7; //] 
    18'h19668: Data = 4'h4; //> 
    18'h19669: Data = 4'h4; //> 
    18'h19670: Data = 4'h4; //> 
    18'h19671: Data = 4'h4; //> 
    18'h19672: Data = 4'ha; //0 
    18'h19673: Data = 4'h2; //+ 
    18'h19674: Data = 4'h4; //> 
    18'h19675: Data = 4'h4; //> 
    18'h19676: Data = 4'h4; //> 
    18'h19677: Data = 4'h4; //> 
    18'h19678: Data = 4'h4; //> 
    18'h19679: Data = 4'h6; //[ 
    18'h19680: Data = 4'h4; //> 
    18'h19681: Data = 4'h4; //> 
    18'h19682: Data = 4'h4; //> 
    18'h19683: Data = 4'h4; //> 
    18'h19684: Data = 4'h4; //> 
    18'h19685: Data = 4'h4; //> 
    18'h19686: Data = 4'h4; //> 
    18'h19687: Data = 4'h4; //> 
    18'h19688: Data = 4'h4; //> 
    18'h19689: Data = 4'h7; //] 
    18'h19690: Data = 4'h4; //> 
    18'h19691: Data = 4'h2; //+ 
    18'h19692: Data = 4'h5; //< 
    18'h19693: Data = 4'h7; //] 
    18'h19694: Data = 4'h7; //] 
    18'h19695: Data = 4'h2; //+ 
    18'h19696: Data = 4'h4; //> 
    18'h19697: Data = 4'h4; //> 
    18'h19698: Data = 4'h4; //> 
    18'h19699: Data = 4'h4; //> 
    18'h19700: Data = 4'h4; //> 
    18'h19701: Data = 4'h4; //> 
    18'h19702: Data = 4'h4; //> 
    18'h19703: Data = 4'h6; //[ 
    18'h19704: Data = 4'h3; //- 
    18'h19705: Data = 4'h5; //< 
    18'h19706: Data = 4'h5; //< 
    18'h19707: Data = 4'h5; //< 
    18'h19708: Data = 4'h5; //< 
    18'h19709: Data = 4'h5; //< 
    18'h19710: Data = 4'h5; //< 
    18'h19711: Data = 4'h5; //< 
    18'h19712: Data = 4'h3; //- 
    18'h19713: Data = 4'h4; //> 
    18'h19714: Data = 4'h4; //> 
    18'h19715: Data = 4'h4; //> 
    18'h19716: Data = 4'h4; //> 
    18'h19717: Data = 4'h4; //> 
    18'h19718: Data = 4'h4; //> 
    18'h19719: Data = 4'h4; //> 
    18'h19720: Data = 4'h7; //] 
    18'h19721: Data = 4'h2; //+ 
    18'h19722: Data = 4'h5; //< 
    18'h19723: Data = 4'h5; //< 
    18'h19724: Data = 4'h5; //< 
    18'h19725: Data = 4'h5; //< 
    18'h19726: Data = 4'h5; //< 
    18'h19727: Data = 4'h5; //< 
    18'h19728: Data = 4'h5; //< 
    18'h19729: Data = 4'h6; //[ 
    18'h19730: Data = 4'h3; //- 
    18'h19731: Data = 4'h4; //> 
    18'h19732: Data = 4'h4; //> 
    18'h19733: Data = 4'h4; //> 
    18'h19734: Data = 4'h4; //> 
    18'h19735: Data = 4'h4; //> 
    18'h19736: Data = 4'h4; //> 
    18'h19737: Data = 4'h4; //> 
    18'h19738: Data = 4'h3; //- 
    18'h19739: Data = 4'h5; //< 
    18'h19740: Data = 4'h5; //< 
    18'h19741: Data = 4'h6; //[ 
    18'h19742: Data = 4'h3; //- 
    18'h19743: Data = 4'h5; //< 
    18'h19744: Data = 4'h5; //< 
    18'h19745: Data = 4'h5; //< 
    18'h19746: Data = 4'h5; //< 
    18'h19747: Data = 4'h5; //< 
    18'h19748: Data = 4'h2; //+ 
    18'h19749: Data = 4'h4; //> 
    18'h19750: Data = 4'h4; //> 
    18'h19751: Data = 4'h4; //> 
    18'h19752: Data = 4'h4; //> 
    18'h19753: Data = 4'h4; //> 
    18'h19754: Data = 4'h7; //] 
    18'h19755: Data = 4'h5; //< 
    18'h19756: Data = 4'h5; //< 
    18'h19757: Data = 4'h5; //< 
    18'h19758: Data = 4'h5; //< 
    18'h19759: Data = 4'h5; //< 
    18'h19760: Data = 4'h6; //[ 
    18'h19761: Data = 4'h3; //- 
    18'h19762: Data = 4'h4; //> 
    18'h19763: Data = 4'h4; //> 
    18'h19764: Data = 4'h4; //> 
    18'h19765: Data = 4'h4; //> 
    18'h19766: Data = 4'h4; //> 
    18'h19767: Data = 4'h2; //+ 
    18'h19768: Data = 4'h5; //< 
    18'h19769: Data = 4'h5; //< 
    18'h19770: Data = 4'h5; //< 
    18'h19771: Data = 4'h5; //< 
    18'h19772: Data = 4'h5; //< 
    18'h19773: Data = 4'h5; //< 
    18'h19774: Data = 4'h5; //< 
    18'h19775: Data = 4'h5; //< 
    18'h19776: Data = 4'h5; //< 
    18'h19777: Data = 4'h5; //< 
    18'h19778: Data = 4'h5; //< 
    18'h19779: Data = 4'h5; //< 
    18'h19780: Data = 4'h5; //< 
    18'h19781: Data = 4'h5; //< 
    18'h19782: Data = 4'h6; //[ 
    18'h19783: Data = 4'h5; //< 
    18'h19784: Data = 4'h5; //< 
    18'h19785: Data = 4'h5; //< 
    18'h19786: Data = 4'h5; //< 
    18'h19787: Data = 4'h5; //< 
    18'h19788: Data = 4'h5; //< 
    18'h19789: Data = 4'h5; //< 
    18'h19790: Data = 4'h5; //< 
    18'h19791: Data = 4'h5; //< 
    18'h19792: Data = 4'h7; //] 
    18'h19793: Data = 4'h4; //> 
    18'h19794: Data = 4'h4; //> 
    18'h19795: Data = 4'h4; //> 
    18'h19796: Data = 4'ha; //0 
    18'h19797: Data = 4'h2; //+ 
    18'h19798: Data = 4'h4; //> 
    18'h19799: Data = 4'h4; //> 
    18'h19800: Data = 4'h4; //> 
    18'h19801: Data = 4'h4; //> 
    18'h19802: Data = 4'h4; //> 
    18'h19803: Data = 4'h4; //> 
    18'h19804: Data = 4'h6; //[ 
    18'h19805: Data = 4'h4; //> 
    18'h19806: Data = 4'h4; //> 
    18'h19807: Data = 4'h4; //> 
    18'h19808: Data = 4'h4; //> 
    18'h19809: Data = 4'h4; //> 
    18'h19810: Data = 4'h4; //> 
    18'h19811: Data = 4'h4; //> 
    18'h19812: Data = 4'h4; //> 
    18'h19813: Data = 4'h4; //> 
    18'h19814: Data = 4'h7; //] 
    18'h19815: Data = 4'h4; //> 
    18'h19816: Data = 4'ha; //0 
    18'h19817: Data = 4'h2; //+ 
    18'h19818: Data = 4'h5; //< 
    18'h19819: Data = 4'h7; //] 
    18'h19820: Data = 4'h7; //] 
    18'h19821: Data = 4'h2; //+ 
    18'h19822: Data = 4'h4; //> 
    18'h19823: Data = 4'h6; //[ 
    18'h19824: Data = 4'h3; //- 
    18'h19825: Data = 4'h5; //< 
    18'h19826: Data = 4'h6; //[ 
    18'h19827: Data = 4'h4; //> 
    18'h19828: Data = 4'h4; //> 
    18'h19829: Data = 4'h4; //> 
    18'h19830: Data = 4'h4; //> 
    18'h19831: Data = 4'h4; //> 
    18'h19832: Data = 4'h4; //> 
    18'h19833: Data = 4'h4; //> 
    18'h19834: Data = 4'h4; //> 
    18'h19835: Data = 4'h4; //> 
    18'h19836: Data = 4'h7; //] 
    18'h19837: Data = 4'h5; //< 
    18'h19838: Data = 4'h5; //< 
    18'h19839: Data = 4'h5; //< 
    18'h19840: Data = 4'h5; //< 
    18'h19841: Data = 4'h5; //< 
    18'h19842: Data = 4'h5; //< 
    18'h19843: Data = 4'h5; //< 
    18'h19844: Data = 4'h5; //< 
    18'h19845: Data = 4'h7; //] 
    18'h19846: Data = 4'h4; //> 
    18'h19847: Data = 4'h4; //> 
    18'h19848: Data = 4'h4; //> 
    18'h19849: Data = 4'h4; //> 
    18'h19850: Data = 4'h4; //> 
    18'h19851: Data = 4'h4; //> 
    18'h19852: Data = 4'h4; //> 
    18'h19853: Data = 4'h4; //> 
    18'h19854: Data = 4'h7; //] 
    18'h19855: Data = 4'h5; //< 
    18'h19856: Data = 4'h5; //< 
    18'h19857: Data = 4'h5; //< 
    18'h19858: Data = 4'h5; //< 
    18'h19859: Data = 4'h5; //< 
    18'h19860: Data = 4'h5; //< 
    18'h19861: Data = 4'h5; //< 
    18'h19862: Data = 4'h5; //< 
    18'h19863: Data = 4'h5; //< 
    18'h19864: Data = 4'h6; //[ 
    18'h19865: Data = 4'h5; //< 
    18'h19866: Data = 4'h5; //< 
    18'h19867: Data = 4'h5; //< 
    18'h19868: Data = 4'h5; //< 
    18'h19869: Data = 4'h5; //< 
    18'h19870: Data = 4'h5; //< 
    18'h19871: Data = 4'h5; //< 
    18'h19872: Data = 4'h5; //< 
    18'h19873: Data = 4'h5; //< 
    18'h19874: Data = 4'h7; //] 
    18'h19875: Data = 4'h4; //> 
    18'h19876: Data = 4'h4; //> 
    18'h19877: Data = 4'h4; //> 
    18'h19878: Data = 4'h4; //> 
    18'h19879: Data = 4'ha; //0 
    18'h19880: Data = 4'h5; //< 
    18'h19881: Data = 4'h5; //< 
    18'h19882: Data = 4'h5; //< 
    18'h19883: Data = 4'h2; //+ 
    18'h19884: Data = 4'h2; //+ 
    18'h19885: Data = 4'h2; //+ 
    18'h19886: Data = 4'h2; //+ 
    18'h19887: Data = 4'h2; //+ 
    18'h19888: Data = 4'h6; //[ 
    18'h19889: Data = 4'h3; //- 
    18'h19890: Data = 4'h6; //[ 
    18'h19891: Data = 4'h3; //- 
    18'h19892: Data = 4'h4; //> 
    18'h19893: Data = 4'h4; //> 
    18'h19894: Data = 4'h4; //> 
    18'h19895: Data = 4'h4; //> 
    18'h19896: Data = 4'h4; //> 
    18'h19897: Data = 4'h4; //> 
    18'h19898: Data = 4'h4; //> 
    18'h19899: Data = 4'h4; //> 
    18'h19900: Data = 4'h4; //> 
    18'h19901: Data = 4'h2; //+ 
    18'h19902: Data = 4'h5; //< 
    18'h19903: Data = 4'h5; //< 
    18'h19904: Data = 4'h5; //< 
    18'h19905: Data = 4'h5; //< 
    18'h19906: Data = 4'h5; //< 
    18'h19907: Data = 4'h5; //< 
    18'h19908: Data = 4'h5; //< 
    18'h19909: Data = 4'h5; //< 
    18'h19910: Data = 4'h5; //< 
    18'h19911: Data = 4'h7; //] 
    18'h19912: Data = 4'h4; //> 
    18'h19913: Data = 4'h4; //> 
    18'h19914: Data = 4'h4; //> 
    18'h19915: Data = 4'h4; //> 
    18'h19916: Data = 4'h4; //> 
    18'h19917: Data = 4'h4; //> 
    18'h19918: Data = 4'h4; //> 
    18'h19919: Data = 4'h4; //> 
    18'h19920: Data = 4'h4; //> 
    18'h19921: Data = 4'h7; //] 
    18'h19922: Data = 4'h4; //> 
    18'h19923: Data = 4'h4; //> 
    18'h19924: Data = 4'h4; //> 
    18'h19925: Data = 4'h4; //> 
    18'h19926: Data = 4'h3; //- 
    18'h19927: Data = 4'h5; //< 
    18'h19928: Data = 4'h5; //< 
    18'h19929: Data = 4'h5; //< 
    18'h19930: Data = 4'h5; //< 
    18'h19931: Data = 4'h5; //< 
    18'h19932: Data = 4'h6; //[ 
    18'h19933: Data = 4'h5; //< 
    18'h19934: Data = 4'h5; //< 
    18'h19935: Data = 4'h5; //< 
    18'h19936: Data = 4'h5; //< 
    18'h19937: Data = 4'h5; //< 
    18'h19938: Data = 4'h5; //< 
    18'h19939: Data = 4'h5; //< 
    18'h19940: Data = 4'h5; //< 
    18'h19941: Data = 4'h5; //< 
    18'h19942: Data = 4'h7; //] 
    18'h19943: Data = 4'h7; //] 
    18'h19944: Data = 4'h4; //> 
    18'h19945: Data = 4'h4; //> 
    18'h19946: Data = 4'h4; //> 
    18'h19947: Data = 4'h7; //] 
    18'h19948: Data = 4'h5; //< 
    18'h19949: Data = 4'h5; //< 
    18'h19950: Data = 4'h5; //< 
    18'h19951: Data = 4'h5; //< 
    18'h19952: Data = 4'h8; //. 
    18'h19953: Data = 4'h4; //> 
    18'h19954: Data = 4'h4; //> 
    18'h19955: Data = 4'h4; //> 
    18'h19956: Data = 4'h4; //> 
    18'h19957: Data = 4'h4; //> 
    18'h19958: Data = 4'h4; //> 
    18'h19959: Data = 4'h4; //> 
    18'h19960: Data = 4'h4; //> 
    18'h19961: Data = 4'h4; //> 
    18'h19962: Data = 4'h4; //> 
    18'h19963: Data = 4'h6; //[ 
    18'h19964: Data = 4'h4; //> 
    18'h19965: Data = 4'h4; //> 
    18'h19966: Data = 4'h4; //> 
    18'h19967: Data = 4'h4; //> 
    18'h19968: Data = 4'h4; //> 
    18'h19969: Data = 4'h4; //> 
    18'h19970: Data = 4'ha; //0 
    18'h19971: Data = 4'h4; //> 
    18'h19972: Data = 4'h4; //> 
    18'h19973: Data = 4'h4; //> 
    18'h19974: Data = 4'h7; //] 
    18'h19975: Data = 4'h5; //< 
    18'h19976: Data = 4'h5; //< 
    18'h19977: Data = 4'h5; //< 
    18'h19978: Data = 4'h5; //< 
    18'h19979: Data = 4'h5; //< 
    18'h19980: Data = 4'h5; //< 
    18'h19981: Data = 4'h5; //< 
    18'h19982: Data = 4'h5; //< 
    18'h19983: Data = 4'h5; //< 
    18'h19984: Data = 4'h6; //[ 
    18'h19985: Data = 4'h5; //< 
    18'h19986: Data = 4'h5; //< 
    18'h19987: Data = 4'h5; //< 
    18'h19988: Data = 4'h5; //< 
    18'h19989: Data = 4'h5; //< 
    18'h19990: Data = 4'h5; //< 
    18'h19991: Data = 4'h5; //< 
    18'h19992: Data = 4'h5; //< 
    18'h19993: Data = 4'h5; //< 
    18'h19994: Data = 4'h7; //] 
    18'h19995: Data = 4'h4; //> 
    18'h19996: Data = 4'h2; //+ 
    18'h19997: Data = 4'h2; //+ 
    18'h19998: Data = 4'h2; //+ 
    18'h19999: Data = 4'h2; //+ 
    18'h20000: Data = 4'h2; //+ 
    18'h20001: Data = 4'h2; //+ 
    18'h20002: Data = 4'h2; //+ 
    18'h20003: Data = 4'h2; //+ 
    18'h20004: Data = 4'h2; //+ 
    18'h20005: Data = 4'h2; //+ 
    18'h20006: Data = 4'h6; //[ 
    18'h20007: Data = 4'h3; //- 
    18'h20008: Data = 4'h6; //[ 
    18'h20009: Data = 4'h3; //- 
    18'h20010: Data = 4'h4; //> 
    18'h20011: Data = 4'h4; //> 
    18'h20012: Data = 4'h4; //> 
    18'h20013: Data = 4'h4; //> 
    18'h20014: Data = 4'h4; //> 
    18'h20015: Data = 4'h4; //> 
    18'h20016: Data = 4'h4; //> 
    18'h20017: Data = 4'h4; //> 
    18'h20018: Data = 4'h4; //> 
    18'h20019: Data = 4'h2; //+ 
    18'h20020: Data = 4'h5; //< 
    18'h20021: Data = 4'h5; //< 
    18'h20022: Data = 4'h5; //< 
    18'h20023: Data = 4'h5; //< 
    18'h20024: Data = 4'h5; //< 
    18'h20025: Data = 4'h5; //< 
    18'h20026: Data = 4'h5; //< 
    18'h20027: Data = 4'h5; //< 
    18'h20028: Data = 4'h5; //< 
    18'h20029: Data = 4'h7; //] 
    18'h20030: Data = 4'h4; //> 
    18'h20031: Data = 4'h4; //> 
    18'h20032: Data = 4'h4; //> 
    18'h20033: Data = 4'h4; //> 
    18'h20034: Data = 4'h4; //> 
    18'h20035: Data = 4'h4; //> 
    18'h20036: Data = 4'h4; //> 
    18'h20037: Data = 4'h4; //> 
    18'h20038: Data = 4'h4; //> 
    18'h20039: Data = 4'h7; //] 
    18'h20040: Data = 4'h4; //> 
    18'h20041: Data = 4'h4; //> 
    18'h20042: Data = 4'h4; //> 
    18'h20043: Data = 4'h4; //> 
    18'h20044: Data = 4'h4; //> 
    18'h20045: Data = 4'h2; //+ 
    18'h20046: Data = 4'h4; //> 
    18'h20047: Data = 4'h4; //> 
    18'h20048: Data = 4'h4; //> 
    18'h20049: Data = 4'h4; //> 
    18'h20050: Data = 4'h4; //> 
    18'h20051: Data = 4'h4; //> 
    18'h20052: Data = 4'h4; //> 
    18'h20053: Data = 4'h4; //> 
    18'h20054: Data = 4'h4; //> 
    18'h20055: Data = 4'h2; //+ 
    18'h20056: Data = 4'h5; //< 
    18'h20057: Data = 4'h5; //< 
    18'h20058: Data = 4'h5; //< 
    18'h20059: Data = 4'h5; //< 
    18'h20060: Data = 4'h5; //< 
    18'h20061: Data = 4'h5; //< 
    18'h20062: Data = 4'h5; //< 
    18'h20063: Data = 4'h5; //< 
    18'h20064: Data = 4'h5; //< 
    18'h20065: Data = 4'h5; //< 
    18'h20066: Data = 4'h5; //< 
    18'h20067: Data = 4'h5; //< 
    18'h20068: Data = 4'h5; //< 
    18'h20069: Data = 4'h5; //< 
    18'h20070: Data = 4'h5; //< 
    18'h20071: Data = 4'h6; //[ 
    18'h20072: Data = 4'h5; //< 
    18'h20073: Data = 4'h5; //< 
    18'h20074: Data = 4'h5; //< 
    18'h20075: Data = 4'h5; //< 
    18'h20076: Data = 4'h5; //< 
    18'h20077: Data = 4'h5; //< 
    18'h20078: Data = 4'h5; //< 
    18'h20079: Data = 4'h5; //< 
    18'h20080: Data = 4'h5; //< 
    18'h20081: Data = 4'h7; //] 
    18'h20082: Data = 4'h4; //> 
    18'h20083: Data = 4'h4; //> 
    18'h20084: Data = 4'h4; //> 
    18'h20085: Data = 4'h4; //> 
    18'h20086: Data = 4'h4; //> 
    18'h20087: Data = 4'h4; //> 
    18'h20088: Data = 4'h4; //> 
    18'h20089: Data = 4'h4; //> 
    18'h20090: Data = 4'h6; //[ 
    18'h20091: Data = 4'h3; //- 
    18'h20092: Data = 4'h5; //< 
    18'h20093: Data = 4'h5; //< 
    18'h20094: Data = 4'h5; //< 
    18'h20095: Data = 4'h5; //< 
    18'h20096: Data = 4'h5; //< 
    18'h20097: Data = 4'h5; //< 
    18'h20098: Data = 4'h5; //< 
    18'h20099: Data = 4'h5; //< 
    18'h20100: Data = 4'h2; //+ 
    18'h20101: Data = 4'h4; //> 
    18'h20102: Data = 4'h4; //> 
    18'h20103: Data = 4'h4; //> 
    18'h20104: Data = 4'h4; //> 
    18'h20105: Data = 4'h4; //> 
    18'h20106: Data = 4'h4; //> 
    18'h20107: Data = 4'h4; //> 
    18'h20108: Data = 4'h4; //> 
    18'h20109: Data = 4'h7; //] 
    18'h20110: Data = 4'h5; //< 
    18'h20111: Data = 4'h5; //< 
    18'h20112: Data = 4'h5; //< 
    18'h20113: Data = 4'h5; //< 
    18'h20114: Data = 4'h5; //< 
    18'h20115: Data = 4'h5; //< 
    18'h20116: Data = 4'h5; //< 
    18'h20117: Data = 4'h5; //< 
    18'h20118: Data = 4'h6; //[ 
    18'h20119: Data = 4'h3; //- 
    18'h20120: Data = 4'h4; //> 
    18'h20121: Data = 4'h4; //> 
    18'h20122: Data = 4'h4; //> 
    18'h20123: Data = 4'h4; //> 
    18'h20124: Data = 4'h4; //> 
    18'h20125: Data = 4'h4; //> 
    18'h20126: Data = 4'h4; //> 
    18'h20127: Data = 4'h4; //> 
    18'h20128: Data = 4'h2; //+ 
    18'h20129: Data = 4'ha; //0 
    18'h20130: Data = 4'h4; //> 
    18'h20131: Data = 4'h6; //[ 
    18'h20132: Data = 4'h4; //> 
    18'h20133: Data = 4'h4; //> 
    18'h20134: Data = 4'h4; //> 
    18'h20135: Data = 4'h4; //> 
    18'h20136: Data = 4'h4; //> 
    18'h20137: Data = 4'h4; //> 
    18'h20138: Data = 4'h4; //> 
    18'h20139: Data = 4'h4; //> 
    18'h20140: Data = 4'h4; //> 
    18'h20141: Data = 4'h7; //] 
    18'h20142: Data = 4'h5; //< 
    18'h20143: Data = 4'h5; //< 
    18'h20144: Data = 4'h5; //< 
    18'h20145: Data = 4'h5; //< 
    18'h20146: Data = 4'h5; //< 
    18'h20147: Data = 4'h5; //< 
    18'h20148: Data = 4'h5; //< 
    18'h20149: Data = 4'h5; //< 
    18'h20150: Data = 4'h5; //< 
    18'h20151: Data = 4'h6; //[ 
    18'h20152: Data = 4'h4; //> 
    18'h20153: Data = 4'h4; //> 
    18'h20154: Data = 4'h4; //> 
    18'h20155: Data = 4'h4; //> 
    18'h20156: Data = 4'h4; //> 
    18'h20157: Data = 4'h4; //> 
    18'h20158: Data = 4'h4; //> 
    18'h20159: Data = 4'h4; //> 
    18'h20160: Data = 4'h6; //[ 
    18'h20161: Data = 4'h3; //- 
    18'h20162: Data = 4'h5; //< 
    18'h20163: Data = 4'h5; //< 
    18'h20164: Data = 4'h5; //< 
    18'h20165: Data = 4'h5; //< 
    18'h20166: Data = 4'h5; //< 
    18'h20167: Data = 4'h5; //< 
    18'h20168: Data = 4'h5; //< 
    18'h20169: Data = 4'h2; //+ 
    18'h20170: Data = 4'h4; //> 
    18'h20171: Data = 4'h4; //> 
    18'h20172: Data = 4'h4; //> 
    18'h20173: Data = 4'h4; //> 
    18'h20174: Data = 4'h4; //> 
    18'h20175: Data = 4'h4; //> 
    18'h20176: Data = 4'h4; //> 
    18'h20177: Data = 4'h7; //] 
    18'h20178: Data = 4'h5; //< 
    18'h20179: Data = 4'h5; //< 
    18'h20180: Data = 4'h5; //< 
    18'h20181: Data = 4'h5; //< 
    18'h20182: Data = 4'h5; //< 
    18'h20183: Data = 4'h5; //< 
    18'h20184: Data = 4'h5; //< 
    18'h20185: Data = 4'h6; //[ 
    18'h20186: Data = 4'h3; //- 
    18'h20187: Data = 4'h4; //> 
    18'h20188: Data = 4'h4; //> 
    18'h20189: Data = 4'h4; //> 
    18'h20190: Data = 4'h4; //> 
    18'h20191: Data = 4'h4; //> 
    18'h20192: Data = 4'h4; //> 
    18'h20193: Data = 4'h4; //> 
    18'h20194: Data = 4'h2; //+ 
    18'h20195: Data = 4'h5; //< 
    18'h20196: Data = 4'h5; //< 
    18'h20197: Data = 4'h5; //< 
    18'h20198: Data = 4'h5; //< 
    18'h20199: Data = 4'h5; //< 
    18'h20200: Data = 4'h5; //< 
    18'h20201: Data = 4'h5; //< 
    18'h20202: Data = 4'h5; //< 
    18'h20203: Data = 4'h6; //[ 
    18'h20204: Data = 4'h5; //< 
    18'h20205: Data = 4'h5; //< 
    18'h20206: Data = 4'h5; //< 
    18'h20207: Data = 4'h5; //< 
    18'h20208: Data = 4'h5; //< 
    18'h20209: Data = 4'h5; //< 
    18'h20210: Data = 4'h5; //< 
    18'h20211: Data = 4'h5; //< 
    18'h20212: Data = 4'h5; //< 
    18'h20213: Data = 4'h7; //] 
    18'h20214: Data = 4'h4; //> 
    18'h20215: Data = 4'h4; //> 
    18'h20216: Data = 4'h4; //> 
    18'h20217: Data = 4'h4; //> 
    18'h20218: Data = 4'h4; //> 
    18'h20219: Data = 4'h4; //> 
    18'h20220: Data = 4'h4; //> 
    18'h20221: Data = 4'h4; //> 
    18'h20222: Data = 4'ha; //0 
    18'h20223: Data = 4'h2; //+ 
    18'h20224: Data = 4'h4; //> 
    18'h20225: Data = 4'h4; //> 
    18'h20226: Data = 4'h7; //] 
    18'h20227: Data = 4'h5; //< 
    18'h20228: Data = 4'h5; //< 
    18'h20229: Data = 4'h5; //< 
    18'h20230: Data = 4'h5; //< 
    18'h20231: Data = 4'h5; //< 
    18'h20232: Data = 4'h5; //< 
    18'h20233: Data = 4'h5; //< 
    18'h20234: Data = 4'h5; //< 
    18'h20235: Data = 4'h5; //< 
    18'h20236: Data = 4'h5; //< 
    18'h20237: Data = 4'h7; //] 
    18'h20238: Data = 4'h7; //] 
    18'h20239: Data = 4'h4; //> 
    18'h20240: Data = 4'h4; //> 
    18'h20241: Data = 4'h4; //> 
    18'h20242: Data = 4'h4; //> 
    18'h20243: Data = 4'h4; //> 
    18'h20244: Data = 4'h4; //> 
    18'h20245: Data = 4'h4; //> 
    18'h20246: Data = 4'h4; //> 
    18'h20247: Data = 4'h6; //[ 
    18'h20248: Data = 4'h3; //- 
    18'h20249: Data = 4'h5; //< 
    18'h20250: Data = 4'h5; //< 
    18'h20251: Data = 4'h5; //< 
    18'h20252: Data = 4'h5; //< 
    18'h20253: Data = 4'h5; //< 
    18'h20254: Data = 4'h5; //< 
    18'h20255: Data = 4'h5; //< 
    18'h20256: Data = 4'h5; //< 
    18'h20257: Data = 4'h2; //+ 
    18'h20258: Data = 4'h4; //> 
    18'h20259: Data = 4'h4; //> 
    18'h20260: Data = 4'h4; //> 
    18'h20261: Data = 4'h4; //> 
    18'h20262: Data = 4'h4; //> 
    18'h20263: Data = 4'h4; //> 
    18'h20264: Data = 4'h4; //> 
    18'h20265: Data = 4'h4; //> 
    18'h20266: Data = 4'h7; //] 
    18'h20267: Data = 4'h5; //< 
    18'h20268: Data = 4'h5; //< 
    18'h20269: Data = 4'h5; //< 
    18'h20270: Data = 4'h5; //< 
    18'h20271: Data = 4'h5; //< 
    18'h20272: Data = 4'h5; //< 
    18'h20273: Data = 4'h5; //< 
    18'h20274: Data = 4'h5; //< 
    18'h20275: Data = 4'h6; //[ 
    18'h20276: Data = 4'h3; //- 
    18'h20277: Data = 4'h4; //> 
    18'h20278: Data = 4'h4; //> 
    18'h20279: Data = 4'h4; //> 
    18'h20280: Data = 4'h4; //> 
    18'h20281: Data = 4'h4; //> 
    18'h20282: Data = 4'h4; //> 
    18'h20283: Data = 4'h4; //> 
    18'h20284: Data = 4'h4; //> 
    18'h20285: Data = 4'h2; //+ 
    18'h20286: Data = 4'h4; //> 
    18'h20287: Data = 4'h6; //[ 
    18'h20288: Data = 4'h4; //> 
    18'h20289: Data = 4'h2; //+ 
    18'h20290: Data = 4'h4; //> 
    18'h20291: Data = 4'h4; //> 
    18'h20292: Data = 4'h4; //> 
    18'h20293: Data = 4'h4; //> 
    18'h20294: Data = 4'h4; //> 
    18'h20295: Data = 4'h6; //[ 
    18'h20296: Data = 4'h3; //- 
    18'h20297: Data = 4'h5; //< 
    18'h20298: Data = 4'h5; //< 
    18'h20299: Data = 4'h5; //< 
    18'h20300: Data = 4'h5; //< 
    18'h20301: Data = 4'h5; //< 
    18'h20302: Data = 4'h3; //- 
    18'h20303: Data = 4'h4; //> 
    18'h20304: Data = 4'h4; //> 
    18'h20305: Data = 4'h4; //> 
    18'h20306: Data = 4'h4; //> 
    18'h20307: Data = 4'h4; //> 
    18'h20308: Data = 4'h7; //] 
    18'h20309: Data = 4'h5; //< 
    18'h20310: Data = 4'h5; //< 
    18'h20311: Data = 4'h5; //< 
    18'h20312: Data = 4'h5; //< 
    18'h20313: Data = 4'h5; //< 
    18'h20314: Data = 4'h6; //[ 
    18'h20315: Data = 4'h3; //- 
    18'h20316: Data = 4'h4; //> 
    18'h20317: Data = 4'h4; //> 
    18'h20318: Data = 4'h4; //> 
    18'h20319: Data = 4'h4; //> 
    18'h20320: Data = 4'h4; //> 
    18'h20321: Data = 4'h2; //+ 
    18'h20322: Data = 4'h5; //< 
    18'h20323: Data = 4'h5; //< 
    18'h20324: Data = 4'h5; //< 
    18'h20325: Data = 4'h5; //< 
    18'h20326: Data = 4'h5; //< 
    18'h20327: Data = 4'h7; //] 
    18'h20328: Data = 4'h4; //> 
    18'h20329: Data = 4'h4; //> 
    18'h20330: Data = 4'h4; //> 
    18'h20331: Data = 4'h4; //> 
    18'h20332: Data = 4'h4; //> 
    18'h20333: Data = 4'h4; //> 
    18'h20334: Data = 4'h4; //> 
    18'h20335: Data = 4'h4; //> 
    18'h20336: Data = 4'h7; //] 
    18'h20337: Data = 4'h5; //< 
    18'h20338: Data = 4'h2; //+ 
    18'h20339: Data = 4'h5; //< 
    18'h20340: Data = 4'h5; //< 
    18'h20341: Data = 4'h5; //< 
    18'h20342: Data = 4'h5; //< 
    18'h20343: Data = 4'h5; //< 
    18'h20344: Data = 4'h5; //< 
    18'h20345: Data = 4'h5; //< 
    18'h20346: Data = 4'h5; //< 
    18'h20347: Data = 4'h6; //[ 
    18'h20348: Data = 4'h4; //> 
    18'h20349: Data = 4'h4; //> 
    18'h20350: Data = 4'h4; //> 
    18'h20351: Data = 4'h4; //> 
    18'h20352: Data = 4'h4; //> 
    18'h20353: Data = 4'h4; //> 
    18'h20354: Data = 4'h6; //[ 
    18'h20355: Data = 4'h3; //- 
    18'h20356: Data = 4'h4; //> 
    18'h20357: Data = 4'h4; //> 
    18'h20358: Data = 4'h2; //+ 
    18'h20359: Data = 4'h5; //< 
    18'h20360: Data = 4'h5; //< 
    18'h20361: Data = 4'h7; //] 
    18'h20362: Data = 4'h5; //< 
    18'h20363: Data = 4'h5; //< 
    18'h20364: Data = 4'h5; //< 
    18'h20365: Data = 4'h5; //< 
    18'h20366: Data = 4'h5; //< 
    18'h20367: Data = 4'h5; //< 
    18'h20368: Data = 4'h5; //< 
    18'h20369: Data = 4'h5; //< 
    18'h20370: Data = 4'h5; //< 
    18'h20371: Data = 4'h5; //< 
    18'h20372: Data = 4'h5; //< 
    18'h20373: Data = 4'h5; //< 
    18'h20374: Data = 4'h5; //< 
    18'h20375: Data = 4'h5; //< 
    18'h20376: Data = 4'h5; //< 
    18'h20377: Data = 4'h7; //] 
    18'h20378: Data = 4'h4; //> 
    18'h20379: Data = 4'h4; //> 
    18'h20380: Data = 4'h4; //> 
    18'h20381: Data = 4'h4; //> 
    18'h20382: Data = 4'h4; //> 
    18'h20383: Data = 4'h4; //> 
    18'h20384: Data = 4'h4; //> 
    18'h20385: Data = 4'h4; //> 
    18'h20386: Data = 4'h4; //> 
    18'h20387: Data = 4'h6; //[ 
    18'h20388: Data = 4'h4; //> 
    18'h20389: Data = 4'h4; //> 
    18'h20390: Data = 4'h4; //> 
    18'h20391: Data = 4'h4; //> 
    18'h20392: Data = 4'h4; //> 
    18'h20393: Data = 4'h4; //> 
    18'h20394: Data = 4'h4; //> 
    18'h20395: Data = 4'h4; //> 
    18'h20396: Data = 4'h4; //> 
    18'h20397: Data = 4'h7; //] 
    18'h20398: Data = 4'h5; //< 
    18'h20399: Data = 4'h5; //< 
    18'h20400: Data = 4'h5; //< 
    18'h20401: Data = 4'h5; //< 
    18'h20402: Data = 4'h5; //< 
    18'h20403: Data = 4'h5; //< 
    18'h20404: Data = 4'h5; //< 
    18'h20405: Data = 4'h5; //< 
    18'h20406: Data = 4'h5; //< 
    18'h20407: Data = 4'h6; //[ 
    18'h20408: Data = 4'h4; //> 
    18'h20409: Data = 4'ha; //0 
    18'h20410: Data = 4'h5; //< 
    18'h20411: Data = 4'h3; //- 
    18'h20412: Data = 4'h4; //> 
    18'h20413: Data = 4'h4; //> 
    18'h20414: Data = 4'h4; //> 
    18'h20415: Data = 4'h4; //> 
    18'h20416: Data = 4'h4; //> 
    18'h20417: Data = 4'h4; //> 
    18'h20418: Data = 4'h4; //> 
    18'h20419: Data = 4'h4; //> 
    18'h20420: Data = 4'h6; //[ 
    18'h20421: Data = 4'h3; //- 
    18'h20422: Data = 4'h5; //< 
    18'h20423: Data = 4'h5; //< 
    18'h20424: Data = 4'h5; //< 
    18'h20425: Data = 4'h5; //< 
    18'h20426: Data = 4'h5; //< 
    18'h20427: Data = 4'h5; //< 
    18'h20428: Data = 4'h5; //< 
    18'h20429: Data = 4'h5; //< 
    18'h20430: Data = 4'h2; //+ 
    18'h20431: Data = 4'h4; //> 
    18'h20432: Data = 4'h6; //[ 
    18'h20433: Data = 4'h5; //< 
    18'h20434: Data = 4'h3; //- 
    18'h20435: Data = 4'h4; //> 
    18'h20436: Data = 4'h3; //- 
    18'h20437: Data = 4'h5; //< 
    18'h20438: Data = 4'h5; //< 
    18'h20439: Data = 4'h2; //+ 
    18'h20440: Data = 4'h4; //> 
    18'h20441: Data = 4'h4; //> 
    18'h20442: Data = 4'h7; //] 
    18'h20443: Data = 4'h5; //< 
    18'h20444: Data = 4'h6; //[ 
    18'h20445: Data = 4'h3; //- 
    18'h20446: Data = 4'h4; //> 
    18'h20447: Data = 4'h2; //+ 
    18'h20448: Data = 4'h5; //< 
    18'h20449: Data = 4'h7; //] 
    18'h20450: Data = 4'h4; //> 
    18'h20451: Data = 4'h4; //> 
    18'h20452: Data = 4'h4; //> 
    18'h20453: Data = 4'h4; //> 
    18'h20454: Data = 4'h4; //> 
    18'h20455: Data = 4'h4; //> 
    18'h20456: Data = 4'h4; //> 
    18'h20457: Data = 4'h4; //> 
    18'h20458: Data = 4'h7; //] 
    18'h20459: Data = 4'h5; //< 
    18'h20460: Data = 4'h5; //< 
    18'h20461: Data = 4'h5; //< 
    18'h20462: Data = 4'h5; //< 
    18'h20463: Data = 4'h5; //< 
    18'h20464: Data = 4'h5; //< 
    18'h20465: Data = 4'h5; //< 
    18'h20466: Data = 4'h6; //[ 
    18'h20467: Data = 4'h3; //- 
    18'h20468: Data = 4'h4; //> 
    18'h20469: Data = 4'h4; //> 
    18'h20470: Data = 4'h4; //> 
    18'h20471: Data = 4'h4; //> 
    18'h20472: Data = 4'h4; //> 
    18'h20473: Data = 4'h4; //> 
    18'h20474: Data = 4'h4; //> 
    18'h20475: Data = 4'h2; //+ 
    18'h20476: Data = 4'h5; //< 
    18'h20477: Data = 4'h5; //< 
    18'h20478: Data = 4'h5; //< 
    18'h20479: Data = 4'h5; //< 
    18'h20480: Data = 4'h5; //< 
    18'h20481: Data = 4'h5; //< 
    18'h20482: Data = 4'h5; //< 
    18'h20483: Data = 4'h7; //] 
    18'h20484: Data = 4'h5; //< 
    18'h20485: Data = 4'h2; //+ 
    18'h20486: Data = 4'h5; //< 
    18'h20487: Data = 4'h5; //< 
    18'h20488: Data = 4'h5; //< 
    18'h20489: Data = 4'h5; //< 
    18'h20490: Data = 4'h5; //< 
    18'h20491: Data = 4'h5; //< 
    18'h20492: Data = 4'h5; //< 
    18'h20493: Data = 4'h5; //< 
    18'h20494: Data = 4'h5; //< 
    18'h20495: Data = 4'h7; //] 
    18'h20496: Data = 4'h4; //> 
    18'h20497: Data = 4'h4; //> 
    18'h20498: Data = 4'h4; //> 
    18'h20499: Data = 4'h4; //> 
    18'h20500: Data = 4'h4; //> 
    18'h20501: Data = 4'h4; //> 
    18'h20502: Data = 4'h4; //> 
    18'h20503: Data = 4'h4; //> 
    18'h20504: Data = 4'h3; //- 
    18'h20505: Data = 4'h5; //< 
    18'h20506: Data = 4'h5; //< 
    18'h20507: Data = 4'h5; //< 
    18'h20508: Data = 4'h5; //< 
    18'h20509: Data = 4'h5; //< 
    18'h20510: Data = 4'ha; //0 
    18'h20511: Data = 4'h2; //+ 
    18'h20512: Data = 4'h5; //< 
    18'h20513: Data = 4'h5; //< 
    18'h20514: Data = 4'h5; //< 
    18'h20515: Data = 4'h7; //] 
    18'h20516: Data = 4'h2; //+ 
    18'h20517: Data = 4'h4; //> 
    18'h20518: Data = 4'h4; //> 
    18'h20519: Data = 4'h4; //> 
    18'h20520: Data = 4'h4; //> 
    18'h20521: Data = 4'h4; //> 
    18'h20522: Data = 4'h4; //> 
    18'h20523: Data = 4'h4; //> 
    18'h20524: Data = 4'h4; //> 
    18'h20525: Data = 4'h6; //[ 
    18'h20526: Data = 4'h3; //- 
    18'h20527: Data = 4'h5; //< 
    18'h20528: Data = 4'h5; //< 
    18'h20529: Data = 4'h5; //< 
    18'h20530: Data = 4'h5; //< 
    18'h20531: Data = 4'h5; //< 
    18'h20532: Data = 4'h5; //< 
    18'h20533: Data = 4'h5; //< 
    18'h20534: Data = 4'h5; //< 
    18'h20535: Data = 4'h3; //- 
    18'h20536: Data = 4'h4; //> 
    18'h20537: Data = 4'h4; //> 
    18'h20538: Data = 4'h4; //> 
    18'h20539: Data = 4'h4; //> 
    18'h20540: Data = 4'h4; //> 
    18'h20541: Data = 4'h4; //> 
    18'h20542: Data = 4'h4; //> 
    18'h20543: Data = 4'h4; //> 
    18'h20544: Data = 4'h7; //] 
    18'h20545: Data = 4'h2; //+ 
    18'h20546: Data = 4'h5; //< 
    18'h20547: Data = 4'h5; //< 
    18'h20548: Data = 4'h5; //< 
    18'h20549: Data = 4'h5; //< 
    18'h20550: Data = 4'h5; //< 
    18'h20551: Data = 4'h5; //< 
    18'h20552: Data = 4'h5; //< 
    18'h20553: Data = 4'h5; //< 
    18'h20554: Data = 4'h6; //[ 
    18'h20555: Data = 4'h3; //- 
    18'h20556: Data = 4'h4; //> 
    18'h20557: Data = 4'h4; //> 
    18'h20558: Data = 4'h4; //> 
    18'h20559: Data = 4'h4; //> 
    18'h20560: Data = 4'h4; //> 
    18'h20561: Data = 4'h4; //> 
    18'h20562: Data = 4'h4; //> 
    18'h20563: Data = 4'h4; //> 
    18'h20564: Data = 4'h3; //- 
    18'h20565: Data = 4'h4; //> 
    18'h20566: Data = 4'h6; //[ 
    18'h20567: Data = 4'h4; //> 
    18'h20568: Data = 4'h4; //> 
    18'h20569: Data = 4'h4; //> 
    18'h20570: Data = 4'h4; //> 
    18'h20571: Data = 4'h4; //> 
    18'h20572: Data = 4'h4; //> 
    18'h20573: Data = 4'h6; //[ 
    18'h20574: Data = 4'h3; //- 
    18'h20575: Data = 4'h4; //> 
    18'h20576: Data = 4'h4; //> 
    18'h20577: Data = 4'h2; //+ 
    18'h20578: Data = 4'h5; //< 
    18'h20579: Data = 4'h5; //< 
    18'h20580: Data = 4'h7; //] 
    18'h20581: Data = 4'h4; //> 
    18'h20582: Data = 4'h4; //> 
    18'h20583: Data = 4'h4; //> 
    18'h20584: Data = 4'h7; //] 
    18'h20585: Data = 4'h5; //< 
    18'h20586: Data = 4'h5; //< 
    18'h20587: Data = 4'h5; //< 
    18'h20588: Data = 4'h5; //< 
    18'h20589: Data = 4'h5; //< 
    18'h20590: Data = 4'h5; //< 
    18'h20591: Data = 4'h5; //< 
    18'h20592: Data = 4'h5; //< 
    18'h20593: Data = 4'h5; //< 
    18'h20594: Data = 4'h6; //[ 
    18'h20595: Data = 4'h4; //> 
    18'h20596: Data = 4'ha; //0 
    18'h20597: Data = 4'h5; //< 
    18'h20598: Data = 4'h3; //- 
    18'h20599: Data = 4'h4; //> 
    18'h20600: Data = 4'h4; //> 
    18'h20601: Data = 4'h4; //> 
    18'h20602: Data = 4'h4; //> 
    18'h20603: Data = 4'h4; //> 
    18'h20604: Data = 4'h4; //> 
    18'h20605: Data = 4'h4; //> 
    18'h20606: Data = 4'h4; //> 
    18'h20607: Data = 4'h6; //[ 
    18'h20608: Data = 4'h3; //- 
    18'h20609: Data = 4'h5; //< 
    18'h20610: Data = 4'h5; //< 
    18'h20611: Data = 4'h5; //< 
    18'h20612: Data = 4'h5; //< 
    18'h20613: Data = 4'h5; //< 
    18'h20614: Data = 4'h5; //< 
    18'h20615: Data = 4'h5; //< 
    18'h20616: Data = 4'h5; //< 
    18'h20617: Data = 4'h2; //+ 
    18'h20618: Data = 4'h4; //> 
    18'h20619: Data = 4'h6; //[ 
    18'h20620: Data = 4'h5; //< 
    18'h20621: Data = 4'h3; //- 
    18'h20622: Data = 4'h4; //> 
    18'h20623: Data = 4'h3; //- 
    18'h20624: Data = 4'h5; //< 
    18'h20625: Data = 4'h5; //< 
    18'h20626: Data = 4'h2; //+ 
    18'h20627: Data = 4'h4; //> 
    18'h20628: Data = 4'h4; //> 
    18'h20629: Data = 4'h7; //] 
    18'h20630: Data = 4'h5; //< 
    18'h20631: Data = 4'h6; //[ 
    18'h20632: Data = 4'h3; //- 
    18'h20633: Data = 4'h4; //> 
    18'h20634: Data = 4'h2; //+ 
    18'h20635: Data = 4'h5; //< 
    18'h20636: Data = 4'h7; //] 
    18'h20637: Data = 4'h4; //> 
    18'h20638: Data = 4'h4; //> 
    18'h20639: Data = 4'h4; //> 
    18'h20640: Data = 4'h4; //> 
    18'h20641: Data = 4'h4; //> 
    18'h20642: Data = 4'h4; //> 
    18'h20643: Data = 4'h4; //> 
    18'h20644: Data = 4'h4; //> 
    18'h20645: Data = 4'h7; //] 
    18'h20646: Data = 4'h5; //< 
    18'h20647: Data = 4'h5; //< 
    18'h20648: Data = 4'h5; //< 
    18'h20649: Data = 4'h5; //< 
    18'h20650: Data = 4'h5; //< 
    18'h20651: Data = 4'h5; //< 
    18'h20652: Data = 4'h5; //< 
    18'h20653: Data = 4'h6; //[ 
    18'h20654: Data = 4'h3; //- 
    18'h20655: Data = 4'h4; //> 
    18'h20656: Data = 4'h4; //> 
    18'h20657: Data = 4'h4; //> 
    18'h20658: Data = 4'h4; //> 
    18'h20659: Data = 4'h4; //> 
    18'h20660: Data = 4'h4; //> 
    18'h20661: Data = 4'h4; //> 
    18'h20662: Data = 4'h2; //+ 
    18'h20663: Data = 4'h5; //< 
    18'h20664: Data = 4'h5; //< 
    18'h20665: Data = 4'h5; //< 
    18'h20666: Data = 4'h5; //< 
    18'h20667: Data = 4'h5; //< 
    18'h20668: Data = 4'h5; //< 
    18'h20669: Data = 4'h5; //< 
    18'h20670: Data = 4'h7; //] 
    18'h20671: Data = 4'h5; //< 
    18'h20672: Data = 4'h2; //+ 
    18'h20673: Data = 4'h5; //< 
    18'h20674: Data = 4'h5; //< 
    18'h20675: Data = 4'h5; //< 
    18'h20676: Data = 4'h5; //< 
    18'h20677: Data = 4'h5; //< 
    18'h20678: Data = 4'h5; //< 
    18'h20679: Data = 4'h5; //< 
    18'h20680: Data = 4'h5; //< 
    18'h20681: Data = 4'h5; //< 
    18'h20682: Data = 4'h7; //] 
    18'h20683: Data = 4'h4; //> 
    18'h20684: Data = 4'h2; //+ 
    18'h20685: Data = 4'h2; //+ 
    18'h20686: Data = 4'h2; //+ 
    18'h20687: Data = 4'h2; //+ 
    18'h20688: Data = 4'h2; //+ 
    18'h20689: Data = 4'h6; //[ 
    18'h20690: Data = 4'h3; //- 
    18'h20691: Data = 4'h6; //[ 
    18'h20692: Data = 4'h3; //- 
    18'h20693: Data = 4'h4; //> 
    18'h20694: Data = 4'h4; //> 
    18'h20695: Data = 4'h4; //> 
    18'h20696: Data = 4'h4; //> 
    18'h20697: Data = 4'h4; //> 
    18'h20698: Data = 4'h4; //> 
    18'h20699: Data = 4'h4; //> 
    18'h20700: Data = 4'h4; //> 
    18'h20701: Data = 4'h4; //> 
    18'h20702: Data = 4'h2; //+ 
    18'h20703: Data = 4'h5; //< 
    18'h20704: Data = 4'h5; //< 
    18'h20705: Data = 4'h5; //< 
    18'h20706: Data = 4'h5; //< 
    18'h20707: Data = 4'h5; //< 
    18'h20708: Data = 4'h5; //< 
    18'h20709: Data = 4'h5; //< 
    18'h20710: Data = 4'h5; //< 
    18'h20711: Data = 4'h5; //< 
    18'h20712: Data = 4'h7; //] 
    18'h20713: Data = 4'h4; //> 
    18'h20714: Data = 4'h4; //> 
    18'h20715: Data = 4'h4; //> 
    18'h20716: Data = 4'h4; //> 
    18'h20717: Data = 4'h4; //> 
    18'h20718: Data = 4'h4; //> 
    18'h20719: Data = 4'h4; //> 
    18'h20720: Data = 4'h4; //> 
    18'h20721: Data = 4'h4; //> 
    18'h20722: Data = 4'h7; //] 
    18'h20723: Data = 4'h4; //> 
    18'h20724: Data = 4'h4; //> 
    18'h20725: Data = 4'h4; //> 
    18'h20726: Data = 4'h4; //> 
    18'h20727: Data = 4'h4; //> 
    18'h20728: Data = 4'h2; //+ 
    18'h20729: Data = 4'h4; //> 
    18'h20730: Data = 4'h4; //> 
    18'h20731: Data = 4'h4; //> 
    18'h20732: Data = 4'h4; //> 
    18'h20733: Data = 4'h4; //> 
    18'h20734: Data = 4'h4; //> 
    18'h20735: Data = 4'h4; //> 
    18'h20736: Data = 4'h4; //> 
    18'h20737: Data = 4'h4; //> 
    18'h20738: Data = 4'h4; //> 
    18'h20739: Data = 4'h4; //> 
    18'h20740: Data = 4'h4; //> 
    18'h20741: Data = 4'h4; //> 
    18'h20742: Data = 4'h4; //> 
    18'h20743: Data = 4'h4; //> 
    18'h20744: Data = 4'h4; //> 
    18'h20745: Data = 4'h4; //> 
    18'h20746: Data = 4'h4; //> 
    18'h20747: Data = 4'h4; //> 
    18'h20748: Data = 4'h4; //> 
    18'h20749: Data = 4'h4; //> 
    18'h20750: Data = 4'h4; //> 
    18'h20751: Data = 4'h4; //> 
    18'h20752: Data = 4'h4; //> 
    18'h20753: Data = 4'h4; //> 
    18'h20754: Data = 4'h4; //> 
    18'h20755: Data = 4'h4; //> 
    18'h20756: Data = 4'h2; //+ 
    18'h20757: Data = 4'h5; //< 
    18'h20758: Data = 4'h5; //< 
    18'h20759: Data = 4'h5; //< 
    18'h20760: Data = 4'h5; //< 
    18'h20761: Data = 4'h5; //< 
    18'h20762: Data = 4'h5; //< 
    18'h20763: Data = 4'h6; //[ 
    18'h20764: Data = 4'h5; //< 
    18'h20765: Data = 4'h5; //< 
    18'h20766: Data = 4'h5; //< 
    18'h20767: Data = 4'h5; //< 
    18'h20768: Data = 4'h5; //< 
    18'h20769: Data = 4'h5; //< 
    18'h20770: Data = 4'h5; //< 
    18'h20771: Data = 4'h5; //< 
    18'h20772: Data = 4'h5; //< 
    18'h20773: Data = 4'h7; //] 
    18'h20774: Data = 4'h4; //> 
    18'h20775: Data = 4'h4; //> 
    18'h20776: Data = 4'h4; //> 
    18'h20777: Data = 4'h4; //> 
    18'h20778: Data = 4'h4; //> 
    18'h20779: Data = 4'h4; //> 
    18'h20780: Data = 4'h4; //> 
    18'h20781: Data = 4'h4; //> 
    18'h20782: Data = 4'h4; //> 
    18'h20783: Data = 4'h6; //[ 
    18'h20784: Data = 4'h4; //> 
    18'h20785: Data = 4'h4; //> 
    18'h20786: Data = 4'h4; //> 
    18'h20787: Data = 4'h4; //> 
    18'h20788: Data = 4'h4; //> 
    18'h20789: Data = 4'h4; //> 
    18'h20790: Data = 4'h6; //[ 
    18'h20791: Data = 4'h3; //- 
    18'h20792: Data = 4'h5; //< 
    18'h20793: Data = 4'h5; //< 
    18'h20794: Data = 4'h5; //< 
    18'h20795: Data = 4'h5; //< 
    18'h20796: Data = 4'h5; //< 
    18'h20797: Data = 4'h5; //< 
    18'h20798: Data = 4'h3; //- 
    18'h20799: Data = 4'h4; //> 
    18'h20800: Data = 4'h4; //> 
    18'h20801: Data = 4'h4; //> 
    18'h20802: Data = 4'h4; //> 
    18'h20803: Data = 4'h4; //> 
    18'h20804: Data = 4'h4; //> 
    18'h20805: Data = 4'h7; //] 
    18'h20806: Data = 4'h2; //+ 
    18'h20807: Data = 4'h5; //< 
    18'h20808: Data = 4'h5; //< 
    18'h20809: Data = 4'h5; //< 
    18'h20810: Data = 4'h5; //< 
    18'h20811: Data = 4'h5; //< 
    18'h20812: Data = 4'h5; //< 
    18'h20813: Data = 4'h6; //[ 
    18'h20814: Data = 4'h3; //- 
    18'h20815: Data = 4'h4; //> 
    18'h20816: Data = 4'h4; //> 
    18'h20817: Data = 4'h4; //> 
    18'h20818: Data = 4'h4; //> 
    18'h20819: Data = 4'h4; //> 
    18'h20820: Data = 4'h4; //> 
    18'h20821: Data = 4'h3; //- 
    18'h20822: Data = 4'h4; //> 
    18'h20823: Data = 4'h4; //> 
    18'h20824: Data = 4'h6; //[ 
    18'h20825: Data = 4'h3; //- 
    18'h20826: Data = 4'h5; //< 
    18'h20827: Data = 4'h5; //< 
    18'h20828: Data = 4'h5; //< 
    18'h20829: Data = 4'h5; //< 
    18'h20830: Data = 4'h5; //< 
    18'h20831: Data = 4'h5; //< 
    18'h20832: Data = 4'h5; //< 
    18'h20833: Data = 4'h5; //< 
    18'h20834: Data = 4'h2; //+ 
    18'h20835: Data = 4'h4; //> 
    18'h20836: Data = 4'h4; //> 
    18'h20837: Data = 4'h4; //> 
    18'h20838: Data = 4'h4; //> 
    18'h20839: Data = 4'h4; //> 
    18'h20840: Data = 4'h4; //> 
    18'h20841: Data = 4'h4; //> 
    18'h20842: Data = 4'h4; //> 
    18'h20843: Data = 4'h7; //] 
    18'h20844: Data = 4'h5; //< 
    18'h20845: Data = 4'h5; //< 
    18'h20846: Data = 4'h5; //< 
    18'h20847: Data = 4'h5; //< 
    18'h20848: Data = 4'h5; //< 
    18'h20849: Data = 4'h5; //< 
    18'h20850: Data = 4'h5; //< 
    18'h20851: Data = 4'h5; //< 
    18'h20852: Data = 4'h6; //[ 
    18'h20853: Data = 4'h3; //- 
    18'h20854: Data = 4'h4; //> 
    18'h20855: Data = 4'h4; //> 
    18'h20856: Data = 4'h4; //> 
    18'h20857: Data = 4'h4; //> 
    18'h20858: Data = 4'h4; //> 
    18'h20859: Data = 4'h4; //> 
    18'h20860: Data = 4'h4; //> 
    18'h20861: Data = 4'h4; //> 
    18'h20862: Data = 4'h2; //+ 
    18'h20863: Data = 4'h5; //< 
    18'h20864: Data = 4'h5; //< 
    18'h20865: Data = 4'h5; //< 
    18'h20866: Data = 4'h5; //< 
    18'h20867: Data = 4'h5; //< 
    18'h20868: Data = 4'h5; //< 
    18'h20869: Data = 4'h5; //< 
    18'h20870: Data = 4'h5; //< 
    18'h20871: Data = 4'h5; //< 
    18'h20872: Data = 4'h5; //< 
    18'h20873: Data = 4'h5; //< 
    18'h20874: Data = 4'h5; //< 
    18'h20875: Data = 4'h5; //< 
    18'h20876: Data = 4'h5; //< 
    18'h20877: Data = 4'h5; //< 
    18'h20878: Data = 4'h5; //< 
    18'h20879: Data = 4'h5; //< 
    18'h20880: Data = 4'h6; //[ 
    18'h20881: Data = 4'h5; //< 
    18'h20882: Data = 4'h5; //< 
    18'h20883: Data = 4'h5; //< 
    18'h20884: Data = 4'h5; //< 
    18'h20885: Data = 4'h5; //< 
    18'h20886: Data = 4'h5; //< 
    18'h20887: Data = 4'h5; //< 
    18'h20888: Data = 4'h5; //< 
    18'h20889: Data = 4'h5; //< 
    18'h20890: Data = 4'h7; //] 
    18'h20891: Data = 4'h4; //> 
    18'h20892: Data = 4'h4; //> 
    18'h20893: Data = 4'h4; //> 
    18'h20894: Data = 4'h4; //> 
    18'h20895: Data = 4'ha; //0 
    18'h20896: Data = 4'h2; //+ 
    18'h20897: Data = 4'h4; //> 
    18'h20898: Data = 4'h4; //> 
    18'h20899: Data = 4'h4; //> 
    18'h20900: Data = 4'h4; //> 
    18'h20901: Data = 4'h4; //> 
    18'h20902: Data = 4'h6; //[ 
    18'h20903: Data = 4'h4; //> 
    18'h20904: Data = 4'h4; //> 
    18'h20905: Data = 4'h4; //> 
    18'h20906: Data = 4'h4; //> 
    18'h20907: Data = 4'h4; //> 
    18'h20908: Data = 4'h4; //> 
    18'h20909: Data = 4'h4; //> 
    18'h20910: Data = 4'h4; //> 
    18'h20911: Data = 4'h4; //> 
    18'h20912: Data = 4'h7; //] 
    18'h20913: Data = 4'h4; //> 
    18'h20914: Data = 4'h2; //+ 
    18'h20915: Data = 4'h5; //< 
    18'h20916: Data = 4'h7; //] 
    18'h20917: Data = 4'h7; //] 
    18'h20918: Data = 4'h2; //+ 
    18'h20919: Data = 4'h4; //> 
    18'h20920: Data = 4'h4; //> 
    18'h20921: Data = 4'h4; //> 
    18'h20922: Data = 4'h4; //> 
    18'h20923: Data = 4'h4; //> 
    18'h20924: Data = 4'h4; //> 
    18'h20925: Data = 4'h4; //> 
    18'h20926: Data = 4'h4; //> 
    18'h20927: Data = 4'h6; //[ 
    18'h20928: Data = 4'h3; //- 
    18'h20929: Data = 4'h5; //< 
    18'h20930: Data = 4'h5; //< 
    18'h20931: Data = 4'h5; //< 
    18'h20932: Data = 4'h5; //< 
    18'h20933: Data = 4'h5; //< 
    18'h20934: Data = 4'h5; //< 
    18'h20935: Data = 4'h5; //< 
    18'h20936: Data = 4'h5; //< 
    18'h20937: Data = 4'h3; //- 
    18'h20938: Data = 4'h4; //> 
    18'h20939: Data = 4'h4; //> 
    18'h20940: Data = 4'h4; //> 
    18'h20941: Data = 4'h4; //> 
    18'h20942: Data = 4'h4; //> 
    18'h20943: Data = 4'h4; //> 
    18'h20944: Data = 4'h4; //> 
    18'h20945: Data = 4'h4; //> 
    18'h20946: Data = 4'h7; //] 
    18'h20947: Data = 4'h2; //+ 
    18'h20948: Data = 4'h5; //< 
    18'h20949: Data = 4'h5; //< 
    18'h20950: Data = 4'h5; //< 
    18'h20951: Data = 4'h5; //< 
    18'h20952: Data = 4'h5; //< 
    18'h20953: Data = 4'h5; //< 
    18'h20954: Data = 4'h5; //< 
    18'h20955: Data = 4'h5; //< 
    18'h20956: Data = 4'h6; //[ 
    18'h20957: Data = 4'h3; //- 
    18'h20958: Data = 4'h4; //> 
    18'h20959: Data = 4'h4; //> 
    18'h20960: Data = 4'h4; //> 
    18'h20961: Data = 4'h4; //> 
    18'h20962: Data = 4'h4; //> 
    18'h20963: Data = 4'h4; //> 
    18'h20964: Data = 4'h4; //> 
    18'h20965: Data = 4'h4; //> 
    18'h20966: Data = 4'h3; //- 
    18'h20967: Data = 4'h5; //< 
    18'h20968: Data = 4'h5; //< 
    18'h20969: Data = 4'h6; //[ 
    18'h20970: Data = 4'h3; //- 
    18'h20971: Data = 4'h5; //< 
    18'h20972: Data = 4'h5; //< 
    18'h20973: Data = 4'h5; //< 
    18'h20974: Data = 4'h5; //< 
    18'h20975: Data = 4'h5; //< 
    18'h20976: Data = 4'h5; //< 
    18'h20977: Data = 4'h2; //+ 
    18'h20978: Data = 4'h4; //> 
    18'h20979: Data = 4'h4; //> 
    18'h20980: Data = 4'h4; //> 
    18'h20981: Data = 4'h4; //> 
    18'h20982: Data = 4'h4; //> 
    18'h20983: Data = 4'h4; //> 
    18'h20984: Data = 4'h7; //] 
    18'h20985: Data = 4'h5; //< 
    18'h20986: Data = 4'h5; //< 
    18'h20987: Data = 4'h5; //< 
    18'h20988: Data = 4'h5; //< 
    18'h20989: Data = 4'h5; //< 
    18'h20990: Data = 4'h5; //< 
    18'h20991: Data = 4'h6; //[ 
    18'h20992: Data = 4'h3; //- 
    18'h20993: Data = 4'h4; //> 
    18'h20994: Data = 4'h4; //> 
    18'h20995: Data = 4'h4; //> 
    18'h20996: Data = 4'h4; //> 
    18'h20997: Data = 4'h4; //> 
    18'h20998: Data = 4'h4; //> 
    18'h20999: Data = 4'h2; //+ 
    18'h21000: Data = 4'h5; //< 
    18'h21001: Data = 4'h5; //< 
    18'h21002: Data = 4'h5; //< 
    18'h21003: Data = 4'h5; //< 
    18'h21004: Data = 4'h5; //< 
    18'h21005: Data = 4'h5; //< 
    18'h21006: Data = 4'h5; //< 
    18'h21007: Data = 4'h5; //< 
    18'h21008: Data = 4'h5; //< 
    18'h21009: Data = 4'h5; //< 
    18'h21010: Data = 4'h5; //< 
    18'h21011: Data = 4'h5; //< 
    18'h21012: Data = 4'h5; //< 
    18'h21013: Data = 4'h5; //< 
    18'h21014: Data = 4'h5; //< 
    18'h21015: Data = 4'h6; //[ 
    18'h21016: Data = 4'h5; //< 
    18'h21017: Data = 4'h5; //< 
    18'h21018: Data = 4'h5; //< 
    18'h21019: Data = 4'h5; //< 
    18'h21020: Data = 4'h5; //< 
    18'h21021: Data = 4'h5; //< 
    18'h21022: Data = 4'h5; //< 
    18'h21023: Data = 4'h5; //< 
    18'h21024: Data = 4'h5; //< 
    18'h21025: Data = 4'h7; //] 
    18'h21026: Data = 4'h4; //> 
    18'h21027: Data = 4'h4; //> 
    18'h21028: Data = 4'h4; //> 
    18'h21029: Data = 4'ha; //0 
    18'h21030: Data = 4'h2; //+ 
    18'h21031: Data = 4'h4; //> 
    18'h21032: Data = 4'h4; //> 
    18'h21033: Data = 4'h4; //> 
    18'h21034: Data = 4'h4; //> 
    18'h21035: Data = 4'h4; //> 
    18'h21036: Data = 4'h4; //> 
    18'h21037: Data = 4'h6; //[ 
    18'h21038: Data = 4'h4; //> 
    18'h21039: Data = 4'h4; //> 
    18'h21040: Data = 4'h4; //> 
    18'h21041: Data = 4'h4; //> 
    18'h21042: Data = 4'h4; //> 
    18'h21043: Data = 4'h4; //> 
    18'h21044: Data = 4'h4; //> 
    18'h21045: Data = 4'h4; //> 
    18'h21046: Data = 4'h4; //> 
    18'h21047: Data = 4'h7; //] 
    18'h21048: Data = 4'h4; //> 
    18'h21049: Data = 4'ha; //0 
    18'h21050: Data = 4'h2; //+ 
    18'h21051: Data = 4'h5; //< 
    18'h21052: Data = 4'h7; //] 
    18'h21053: Data = 4'h7; //] 
    18'h21054: Data = 4'h2; //+ 
    18'h21055: Data = 4'h4; //> 
    18'h21056: Data = 4'h6; //[ 
    18'h21057: Data = 4'h3; //- 
    18'h21058: Data = 4'h5; //< 
    18'h21059: Data = 4'h6; //[ 
    18'h21060: Data = 4'h4; //> 
    18'h21061: Data = 4'h4; //> 
    18'h21062: Data = 4'h4; //> 
    18'h21063: Data = 4'h4; //> 
    18'h21064: Data = 4'h4; //> 
    18'h21065: Data = 4'h4; //> 
    18'h21066: Data = 4'h4; //> 
    18'h21067: Data = 4'h4; //> 
    18'h21068: Data = 4'h4; //> 
    18'h21069: Data = 4'h7; //] 
    18'h21070: Data = 4'h5; //< 
    18'h21071: Data = 4'h5; //< 
    18'h21072: Data = 4'h5; //< 
    18'h21073: Data = 4'h5; //< 
    18'h21074: Data = 4'h5; //< 
    18'h21075: Data = 4'h5; //< 
    18'h21076: Data = 4'h5; //< 
    18'h21077: Data = 4'h5; //< 
    18'h21078: Data = 4'h7; //] 
    18'h21079: Data = 4'h4; //> 
    18'h21080: Data = 4'h4; //> 
    18'h21081: Data = 4'h4; //> 
    18'h21082: Data = 4'h4; //> 
    18'h21083: Data = 4'h4; //> 
    18'h21084: Data = 4'h4; //> 
    18'h21085: Data = 4'h4; //> 
    18'h21086: Data = 4'h4; //> 
    18'h21087: Data = 4'h7; //] 
    18'h21088: Data = 4'h5; //< 
    18'h21089: Data = 4'h5; //< 
    18'h21090: Data = 4'h5; //< 
    18'h21091: Data = 4'h5; //< 
    18'h21092: Data = 4'h5; //< 
    18'h21093: Data = 4'h5; //< 
    18'h21094: Data = 4'h5; //< 
    18'h21095: Data = 4'h5; //< 
    18'h21096: Data = 4'h5; //< 
    18'h21097: Data = 4'h6; //[ 
    18'h21098: Data = 4'h5; //< 
    18'h21099: Data = 4'h5; //< 
    18'h21100: Data = 4'h5; //< 
    18'h21101: Data = 4'h5; //< 
    18'h21102: Data = 4'h5; //< 
    18'h21103: Data = 4'h5; //< 
    18'h21104: Data = 4'h5; //< 
    18'h21105: Data = 4'h5; //< 
    18'h21106: Data = 4'h5; //< 
    18'h21107: Data = 4'h7; //] 
    18'h21108: Data = 4'h4; //> 
    18'h21109: Data = 4'h4; //> 
    18'h21110: Data = 4'h4; //> 
    18'h21111: Data = 4'h4; //> 
    18'h21112: Data = 4'ha; //0 
    18'h21113: Data = 4'h5; //< 
    18'h21114: Data = 4'h5; //< 
    18'h21115: Data = 4'h5; //< 
    18'h21116: Data = 4'h2; //+ 
    18'h21117: Data = 4'h2; //+ 
    18'h21118: Data = 4'h2; //+ 
    18'h21119: Data = 4'h2; //+ 
    18'h21120: Data = 4'h2; //+ 
    18'h21121: Data = 4'h6; //[ 
    18'h21122: Data = 4'h3; //- 
    18'h21123: Data = 4'h6; //[ 
    18'h21124: Data = 4'h3; //- 
    18'h21125: Data = 4'h4; //> 
    18'h21126: Data = 4'h4; //> 
    18'h21127: Data = 4'h4; //> 
    18'h21128: Data = 4'h4; //> 
    18'h21129: Data = 4'h4; //> 
    18'h21130: Data = 4'h4; //> 
    18'h21131: Data = 4'h4; //> 
    18'h21132: Data = 4'h4; //> 
    18'h21133: Data = 4'h4; //> 
    18'h21134: Data = 4'h2; //+ 
    18'h21135: Data = 4'h5; //< 
    18'h21136: Data = 4'h5; //< 
    18'h21137: Data = 4'h5; //< 
    18'h21138: Data = 4'h5; //< 
    18'h21139: Data = 4'h5; //< 
    18'h21140: Data = 4'h5; //< 
    18'h21141: Data = 4'h5; //< 
    18'h21142: Data = 4'h5; //< 
    18'h21143: Data = 4'h5; //< 
    18'h21144: Data = 4'h7; //] 
    18'h21145: Data = 4'h4; //> 
    18'h21146: Data = 4'h4; //> 
    18'h21147: Data = 4'h4; //> 
    18'h21148: Data = 4'h4; //> 
    18'h21149: Data = 4'h4; //> 
    18'h21150: Data = 4'h4; //> 
    18'h21151: Data = 4'h4; //> 
    18'h21152: Data = 4'h4; //> 
    18'h21153: Data = 4'h4; //> 
    18'h21154: Data = 4'h7; //] 
    18'h21155: Data = 4'h4; //> 
    18'h21156: Data = 4'h4; //> 
    18'h21157: Data = 4'h4; //> 
    18'h21158: Data = 4'h4; //> 
    18'h21159: Data = 4'h4; //> 
    18'h21160: Data = 4'h3; //- 
    18'h21161: Data = 4'h4; //> 
    18'h21162: Data = 4'h4; //> 
    18'h21163: Data = 4'h4; //> 
    18'h21164: Data = 4'h4; //> 
    18'h21165: Data = 4'h4; //> 
    18'h21166: Data = 4'h4; //> 
    18'h21167: Data = 4'h4; //> 
    18'h21168: Data = 4'h4; //> 
    18'h21169: Data = 4'h4; //> 
    18'h21170: Data = 4'h4; //> 
    18'h21171: Data = 4'h4; //> 
    18'h21172: Data = 4'h4; //> 
    18'h21173: Data = 4'h4; //> 
    18'h21174: Data = 4'h4; //> 
    18'h21175: Data = 4'h4; //> 
    18'h21176: Data = 4'h4; //> 
    18'h21177: Data = 4'h4; //> 
    18'h21178: Data = 4'h4; //> 
    18'h21179: Data = 4'h4; //> 
    18'h21180: Data = 4'h4; //> 
    18'h21181: Data = 4'h4; //> 
    18'h21182: Data = 4'h4; //> 
    18'h21183: Data = 4'h4; //> 
    18'h21184: Data = 4'h4; //> 
    18'h21185: Data = 4'h4; //> 
    18'h21186: Data = 4'h4; //> 
    18'h21187: Data = 4'h4; //> 
    18'h21188: Data = 4'h3; //- 
    18'h21189: Data = 4'h5; //< 
    18'h21190: Data = 4'h5; //< 
    18'h21191: Data = 4'h5; //< 
    18'h21192: Data = 4'h5; //< 
    18'h21193: Data = 4'h5; //< 
    18'h21194: Data = 4'h5; //< 
    18'h21195: Data = 4'h6; //[ 
    18'h21196: Data = 4'h5; //< 
    18'h21197: Data = 4'h5; //< 
    18'h21198: Data = 4'h5; //< 
    18'h21199: Data = 4'h5; //< 
    18'h21200: Data = 4'h5; //< 
    18'h21201: Data = 4'h5; //< 
    18'h21202: Data = 4'h5; //< 
    18'h21203: Data = 4'h5; //< 
    18'h21204: Data = 4'h5; //< 
    18'h21205: Data = 4'h7; //] 
    18'h21206: Data = 4'h7; //] 
    18'h21207: Data = 4'h4; //> 
    18'h21208: Data = 4'h4; //> 
    18'h21209: Data = 4'h4; //> 
    18'h21210: Data = 4'h7; //] 
    default: Data = {dataSize{1'b0}};
  endcase

/* verilator lint_on WIDTHEXPAND */
endmodule
