module tb;




endmodule