module DekatronCarrySignal(
    input wire [9:0] In,
    output reg CarryLow,
    output reg CarryHigh
); 
/*This module generates carry signal for full 10-position widh dekatron*/

wire carryLowPin = In[0];
wire noCarryPin = In[1] | In[2] | In[3] | In[4] | In[5] | In[6] | In[7] | In[8];
wire carryHighPin = In[9];

always_latch begin
    CarryLow <= carryLowPin ? 1'b1 : (noCarryPin | carryHighPin) ? 1'b0 : CarryLow;
    CarryHigh <= carryHighPin ? 1'b1 : (noCarryPin | carryLowPin) ? 1'b0 : CarryHigh;
end
 
endmodule


